// REVISION    : $Revision: 1.3 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
tx2048x40
#
(
parameter
TABITS
=
12
)
(
CORETSE_AHBI10
,
CORETSE_AHBl10
,
CORETSE_AHBo10
,
CORETSE_AHBi10
,
CORETSE_AHBOo0
,
CORETSE_AHBIo0
,
CORETSE_AHBlo0
)
;
input
CORETSE_AHBI10
;
input
CORETSE_AHBl10
;
input
CORETSE_AHBo10
;
input
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBi10
;
input
[
39
:
0
]
CORETSE_AHBOo0
;
input
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBIo0
;
output
[
39
:
0
]
CORETSE_AHBlo0
;
reg
[
39
:
0
]
CORETSE_AHBlo0
;
parameter
CORETSE_AHBIoII
=
1
;
parameter
CORETSE_AHBOoOoI
=
1
;
parameter
CORETSE_AHBIoOoI
=
4
;
wire
CORETSE_AHBloOoI
;
reg
[
39
:
0
]
CORETSE_AHBooOoI
[
0
:
(
1
<<
TABITS
)
-
1
]
;
assign
#
CORETSE_AHBOoOoI
CORETSE_AHBloOoI
=
CORETSE_AHBI10
;
always
@
(
posedge
CORETSE_AHBloOoI
)
if
(
~
CORETSE_AHBo10
)
CORETSE_AHBooOoI
[
CORETSE_AHBi10
]
=
CORETSE_AHBOo0
;
always
@
(
posedge
CORETSE_AHBl10
)
CORETSE_AHBlo0
=
#
CORETSE_AHBIoOoI
CORETSE_AHBooOoI
[
CORETSE_AHBIo0
]
;
endmodule
