//                        Proprietary and Confidential                          
//                  Copyright (c) 2013 All Rights Reserved                     
// REVISION    : $Revision: 1.9 $                                                  
module
sib_fifo_top
#
(
parameter
CORETSE_AHBIl10I
=
8
,
parameter
CORETSE_AHBll10I
=
4
,
parameter
CORETSE_AHBol10I
=
0
,
parameter
CORETSE_AHBil10I
=
0
,
parameter
CORETSE_AHBO010I
=
0
,
parameter
CORETSE_AHBI010I
=
1
,
parameter
CORETSE_AHBo1IoI
=
0
)
(
input
CORETSE_AHBo010I,
input
CORETSE_AHBi010I,
input
CORETSE_AHBO110I,
input
CORETSE_AHBI110I,
input
[
CORETSE_AHBIl10I
-
1
:
0
]
CORETSE_AHBl110I,
output
[
CORETSE_AHBIl10I
-
1
:
0
]
CORETSE_AHBo110I,
input
CORETSE_AHBi110I,
input
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBOo10I,
output
CORETSE_AHBIo10I,
output
CORETSE_AHBlo10I,
input
CORETSE_AHBOi10I,
input
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBIi10I,
output
[
CORETSE_AHBll10I
:
0
]
CORETSE_AHBoo10I,
output
[
CORETSE_AHBll10I
:
0
]
CORETSE_AHBio10I,
output
CORETSE_AHBli10I,
output
CORETSE_AHBoi10I
)
;
localparam
CORETSE_AHBO1IoI
=
(
1
<<
CORETSE_AHBll10I
)
;
reg
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBi1IoI
,
CORETSE_AHBOoIoI
,
CORETSE_AHBIoIoI
,
CORETSE_AHBloIoI
;
wire
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBooIoI
,
CORETSE_AHBioIoI
,
CORETSE_AHBOiIoI
,
CORETSE_AHBIiIoI
;
reg
[
CORETSE_AHBll10I
:
0
]
CORETSE_AHBliIoI
,
CORETSE_AHBoiIoI
;
reg
CORETSE_AHBiiIoI
,
CORETSE_AHBOOloI
,
CORETSE_AHBIOloI
,
CORETSE_AHBlOloI
;
wire
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBoOloI
,
CORETSE_AHBiOloI
;
assign
CORETSE_AHBIo10I
=
CORETSE_AHBOOloI
;
assign
CORETSE_AHBli10I
=
CORETSE_AHBlOloI
;
assign
CORETSE_AHBlo10I
=
(
CORETSE_AHBliIoI
>=
CORETSE_AHBOo10I
)
;
assign
CORETSE_AHBoi10I
=
(
CORETSE_AHBoiIoI
<=
CORETSE_AHBIi10I
)
;
assign
CORETSE_AHBoo10I
=
CORETSE_AHBliIoI
;
assign
CORETSE_AHBio10I
=
CORETSE_AHBoiIoI
;
assign
CORETSE_AHBOIloI
=
(
CORETSE_AHBi110I
&
!
CORETSE_AHBOOloI
)
;
always
@
(
*
)
begin
if
(
CORETSE_AHBOIloI
)
CORETSE_AHBi1IoI
=
(
CORETSE_AHBOoIoI
==
CORETSE_AHBO1IoI
-
1
)
?
{
CORETSE_AHBll10I
{
1
'b
0
}
}
:
(
CORETSE_AHBOoIoI
+
{
{
(
CORETSE_AHBll10I
-
1
)
{
1
'b
0
}
}
,
1
'b
1
}
)
;
else
CORETSE_AHBi1IoI
=
CORETSE_AHBOoIoI
;
end
always
@
(
*
)
begin
if
(
CORETSE_AHBOOloI
&
(
CORETSE_AHBOoIoI
==
CORETSE_AHBooIoI
)
)
CORETSE_AHBliIoI
=
CORETSE_AHBO1IoI
;
else
if
(
CORETSE_AHBOoIoI
>=
CORETSE_AHBooIoI
)
CORETSE_AHBliIoI
=
(
CORETSE_AHBOoIoI
-
CORETSE_AHBooIoI
)
;
else
CORETSE_AHBliIoI
=
CORETSE_AHBO1IoI
-
(
CORETSE_AHBooIoI
-
CORETSE_AHBOoIoI
)
;
end
always
@
(
*
)
begin
if
(
(
CORETSE_AHBliIoI
==
CORETSE_AHBO1IoI
-
1
)
&
CORETSE_AHBOIloI
&
!
CORETSE_AHBOOloI
)
CORETSE_AHBiiIoI
=
1
'b
1
;
else
if
(
(
CORETSE_AHBOoIoI
!=
CORETSE_AHBooIoI
)
&
CORETSE_AHBOOloI
)
CORETSE_AHBiiIoI
=
1
'b
0
;
else
CORETSE_AHBiiIoI
=
CORETSE_AHBOOloI
;
end
assign
CORETSE_AHBoOloI
=
CORETSE_AHBIIloI
(
CORETSE_AHBOoIoI
)
;
sib_sync_2flp
#
(
.CORETSE_AHBlIloI
(
CORETSE_AHBll10I
)
,
.CORETSE_AHBoIloI
(
CORETSE_AHBo1IoI
)
)
CORETSE_AHBiIloI
(
.CORETSE_AHBOlloI
(
CORETSE_AHBo010I
)
,
.CORETSE_AHBIlloI
(
CORETSE_AHBO110I
)
,
.CORETSE_AHBllloI
(
CORETSE_AHBi010I
)
,
.CORETSE_AHBolloI
(
CORETSE_AHBI110I
)
,
.CORETSE_AHBilloI
(
CORETSE_AHBoOloI
)
,
.CORETSE_AHBO0loI
(
CORETSE_AHBIiIoI
)
)
;
generate
if
(
CORETSE_AHBI010I
==
1
)
assign
CORETSE_AHBOiIoI
=
CORETSE_AHBI0loI
(
CORETSE_AHBIiIoI
)
;
else
assign
CORETSE_AHBOiIoI
=
CORETSE_AHBOoIoI
;
endgenerate
assign
CORETSE_AHBl0loI
=
(
CORETSE_AHBOi10I
&
!
CORETSE_AHBlOloI
)
;
always
@
(
*
)
begin
if
(
CORETSE_AHBl0loI
)
CORETSE_AHBIoIoI
=
(
CORETSE_AHBloIoI
==
CORETSE_AHBO1IoI
-
1
)
?
{
CORETSE_AHBll10I
{
1
'b
0
}
}
:
(
CORETSE_AHBloIoI
+
{
{
(
CORETSE_AHBll10I
-
1
)
{
1
'b
0
}
}
,
1
'b
1
}
)
;
else
CORETSE_AHBIoIoI
=
CORETSE_AHBloIoI
;
end
always
@
(
*
)
begin
if
(
CORETSE_AHBlOloI
&
(
CORETSE_AHBloIoI
==
CORETSE_AHBOiIoI
)
)
CORETSE_AHBoiIoI
=
{
(
CORETSE_AHBll10I
+
1
)
{
1
'b
0
}
}
;
else
if
(
CORETSE_AHBOiIoI
>
CORETSE_AHBloIoI
)
CORETSE_AHBoiIoI
=
(
CORETSE_AHBOiIoI
-
CORETSE_AHBloIoI
)
;
else
CORETSE_AHBoiIoI
=
CORETSE_AHBO1IoI
-
(
CORETSE_AHBloIoI
-
CORETSE_AHBOiIoI
)
;
end
always
@
(
*
)
begin
if
(
(
CORETSE_AHBloIoI
!=
CORETSE_AHBOiIoI
)
&
CORETSE_AHBlOloI
)
CORETSE_AHBIOloI
=
1
'b
0
;
else
if
(
(
CORETSE_AHBoiIoI
==
{
{
CORETSE_AHBll10I
{
1
'b
0
}
}
,
1
'b
1
}
)
&
CORETSE_AHBl0loI
&
!
CORETSE_AHBlOloI
)
CORETSE_AHBIOloI
=
1
'b
1
;
else
CORETSE_AHBIOloI
=
CORETSE_AHBlOloI
;
end
assign
CORETSE_AHBiOloI
=
CORETSE_AHBIIloI
(
CORETSE_AHBloIoI
)
;
sib_sync_2flp
#
(
.CORETSE_AHBlIloI
(
CORETSE_AHBll10I
)
,
.CORETSE_AHBoIloI
(
CORETSE_AHBo1IoI
)
)
CORETSE_AHBo0loI
(
.CORETSE_AHBOlloI
(
CORETSE_AHBO110I
)
,
.CORETSE_AHBIlloI
(
CORETSE_AHBo010I
)
,
.CORETSE_AHBllloI
(
CORETSE_AHBI110I
)
,
.CORETSE_AHBolloI
(
CORETSE_AHBi010I
)
,
.CORETSE_AHBilloI
(
CORETSE_AHBiOloI
)
,
.CORETSE_AHBO0loI
(
CORETSE_AHBioIoI
)
)
;
generate
if
(
CORETSE_AHBI010I
==
1
)
assign
CORETSE_AHBooIoI
=
CORETSE_AHBI0loI
(
CORETSE_AHBioIoI
)
;
else
assign
CORETSE_AHBooIoI
=
CORETSE_AHBloIoI
;
endgenerate
always
@
(
posedge
CORETSE_AHBo010I
or
negedge
CORETSE_AHBi010I
)
begin
if
(
!
CORETSE_AHBi010I
)
begin
CORETSE_AHBOoIoI
<=
{
CORETSE_AHBll10I
{
1
'b
0
}
}
;
CORETSE_AHBOOloI
<=
1
'b
0
;
end
else
begin
CORETSE_AHBOoIoI
<=
CORETSE_AHBi1IoI
;
CORETSE_AHBOOloI
<=
CORETSE_AHBiiIoI
;
end
end
always
@
(
posedge
CORETSE_AHBO110I
or
negedge
CORETSE_AHBI110I
)
begin
if
(
!
CORETSE_AHBI110I
)
begin
CORETSE_AHBloIoI
<=
{
CORETSE_AHBll10I
{
1
'b
0
}
}
;
CORETSE_AHBlOloI
<=
1
'b
1
;
end
else
begin
CORETSE_AHBloIoI
<=
CORETSE_AHBIoIoI
;
CORETSE_AHBlOloI
<=
CORETSE_AHBIOloI
;
end
end
sib_fifo_mem2p
#
(
.CORETSE_AHBIl10I
(
CORETSE_AHBIl10I
)
,
.CORETSE_AHBol10I
(
CORETSE_AHBol10I
)
,
.CORETSE_AHBil10I
(
CORETSE_AHBil10I
)
,
.CORETSE_AHBO010I
(
CORETSE_AHBO010I
)
,
.CORETSE_AHBll10I
(
CORETSE_AHBll10I
)
)
CORETSE_AHBi0loI
(
.CORETSE_AHBo010I
(
CORETSE_AHBo010I
)
,
.CORETSE_AHBO110I
(
CORETSE_AHBO110I
)
,
.CORETSE_AHBI0IoI
(
CORETSE_AHBOIloI
)
,
.CORETSE_AHBl0IoI
(
CORETSE_AHBl0loI
)
,
.CORETSE_AHBo0IoI
(
CORETSE_AHBOoIoI
)
,
.CORETSE_AHBi0IoI
(
CORETSE_AHBloIoI
)
,
.CORETSE_AHBl110I
(
CORETSE_AHBl110I
)
,
.CORETSE_AHBo110I
(
CORETSE_AHBo110I
)
)
;
function
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBI0loI
;
input
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBO1loI
;
integer
CORETSE_AHBOloI
;
begin
for
(
CORETSE_AHBOloI
=
0
;
CORETSE_AHBOloI
<
CORETSE_AHBll10I
;
CORETSE_AHBOloI
=
CORETSE_AHBOloI
+
1
)
CORETSE_AHBI0loI
[
CORETSE_AHBOloI
]
=
^
(
CORETSE_AHBO1loI
>>
CORETSE_AHBOloI
)
;
end
endfunction
function
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBIIloI
;
input
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBI1loI
;
begin
CORETSE_AHBIIloI
=
(
CORETSE_AHBI1loI
>>
1
)
^
CORETSE_AHBI1loI
;
end
endfunction
endmodule
