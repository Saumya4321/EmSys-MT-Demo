// REVISION    : $Revision: 1.1 $
//              Mentor Proprietary and Confidential
//              Copyright (c) 2000, Mentor Intellectual Property Development
`timescale 1ns/1ns
module
pemstat
(
CORETSE_AHBo1Oi
,
CORETSE_AHBi1Oi
,
CORETSE_AHBl1o
,
CORETSE_AHBo1o
,
CORETSE_AHBlOo1
,
CORETSE_AHBIOo1
,
CORETSE_AHBOoOi
,
CORETSE_AHBIoOi
,
CORETSE_AHBloOi
,
CORETSE_AHBooOi
,
CORETSE_AHBioOi
,
CORETSE_AHBOiOi
,
CORETSE_AHBIiOi
,
CORETSE_AHBliOi
,
CORETSE_AHBoiOi
,
CORETSE_AHBiiOi
,
CORETSE_AHBOOIi
,
CORETSE_AHBIOIi
,
CORETSE_AHBlOIi
,
CORETSE_AHBoOIi
)
;
input
CORETSE_AHBo1Oi
,
CORETSE_AHBi1Oi
;
input
CORETSE_AHBo1o
;
input
[
30
:
0
]
CORETSE_AHBl1o
;
input
CORETSE_AHBIOo1
;
input
[
51
:
0
]
CORETSE_AHBlOo1
;
input
CORETSE_AHBOoOi
,
CORETSE_AHBIoOi
;
input
CORETSE_AHBloOi
;
input
CORETSE_AHBooOi
,
CORETSE_AHBioOi
,
CORETSE_AHBOiOi
,
CORETSE_AHBIiOi
;
input
[
6
:
0
]
CORETSE_AHBliOi
;
input
CORETSE_AHBoiOi
,
CORETSE_AHBiiOi
;
input
[
31
:
0
]
CORETSE_AHBOOIi
;
output
[
31
:
0
]
CORETSE_AHBIOIi
;
output
CORETSE_AHBlOIi
,
CORETSE_AHBoOIi
;
wire
[
15
:
0
]
CORETSE_AHBiOIi
;
wire
[
3
:
0
]
CORETSE_AHBOIIi
;
wire
[
43
:
0
]
CORETSE_AHBIIIi
;
wire
[
43
:
0
]
CORETSE_AHBlIIi
;
wire
[
43
:
0
]
CORETSE_AHBoIIi
;
wire
[
43
:
0
]
CORETSE_AHBiIIi
;
wire
[
43
:
0
]
CORETSE_AHBOlIi
;
wire
[
30
:
0
]
CORETSE_AHBIlIi
,
CORETSE_AHBllIi
,
CORETSE_AHBolIi
,
CORETSE_AHBilIi
,
CORETSE_AHBO0Ii
,
CORETSE_AHBI0Ii
,
CORETSE_AHBl0Ii
,
CORETSE_AHBo0Ii
;
wire
[
30
:
0
]
CORETSE_AHBi0Ii
,
CORETSE_AHBO1Ii
,
CORETSE_AHBI1Ii
,
CORETSE_AHBl1Ii
,
CORETSE_AHBo1Ii
,
CORETSE_AHBi1Ii
,
CORETSE_AHBOoIi
,
CORETSE_AHBIoIi
;
wire
[
30
:
0
]
CORETSE_AHBloIi
,
CORETSE_AHBooIi
,
CORETSE_AHBioIi
,
CORETSE_AHBOiIi
,
CORETSE_AHBIiIi
,
CORETSE_AHBliIi
,
CORETSE_AHBoiIi
,
CORETSE_AHBiiIi
;
wire
[
30
:
0
]
CORETSE_AHBOOli
,
CORETSE_AHBIOli
,
CORETSE_AHBlOli
,
CORETSE_AHBoOli
,
CORETSE_AHBiOli
,
CORETSE_AHBOIli
,
CORETSE_AHBIIli
,
CORETSE_AHBlIli
;
wire
[
30
:
0
]
CORETSE_AHBoIli
,
CORETSE_AHBiIli
,
CORETSE_AHBOlli
,
CORETSE_AHBIlli
,
CORETSE_AHBllli
,
CORETSE_AHBolli
,
CORETSE_AHBilli
,
CORETSE_AHBO0li
;
wire
[
30
:
0
]
CORETSE_AHBI0li
,
CORETSE_AHBl0li
,
CORETSE_AHBo0li
,
CORETSE_AHBi0li
;
pemstat_cntrl
CORETSE_AHBO1li
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBlOo1
(
CORETSE_AHBlOo1
)
,
.CORETSE_AHBIOo1
(
CORETSE_AHBIOo1
)
,
.CORETSE_AHBOoOi
(
CORETSE_AHBOoOi
)
,
.CORETSE_AHBIoOi
(
CORETSE_AHBIoOi
)
,
.CORETSE_AHBloOi
(
CORETSE_AHBloOi
)
,
.CORETSE_AHBOiOi
(
CORETSE_AHBOiOi
)
,
.CORETSE_AHBIiOi
(
CORETSE_AHBIiOi
)
,
.CORETSE_AHBiOIi
(
CORETSE_AHBiOIi
)
,
.CORETSE_AHBOIIi
(
CORETSE_AHBOIIi
)
,
.CORETSE_AHBIIIi
(
CORETSE_AHBIIIi
)
)
;
pemstat_store
CORETSE_AHBI1li
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBiOIi
(
CORETSE_AHBiOIi
)
,
.CORETSE_AHBOIIi
(
CORETSE_AHBOIIi
)
,
.CORETSE_AHBIIIi
(
CORETSE_AHBIIIi
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBOOIi
)
,
.CORETSE_AHBOlIi
(
CORETSE_AHBOlIi
)
,
.CORETSE_AHBIlIi
(
CORETSE_AHBIlIi
)
,
.CORETSE_AHBllIi
(
CORETSE_AHBllIi
)
,
.CORETSE_AHBolIi
(
CORETSE_AHBolIi
)
,
.CORETSE_AHBilIi
(
CORETSE_AHBilIi
)
,
.CORETSE_AHBO0Ii
(
CORETSE_AHBO0Ii
)
,
.CORETSE_AHBI0Ii
(
CORETSE_AHBI0Ii
)
,
.CORETSE_AHBl0Ii
(
CORETSE_AHBl0Ii
)
,
.CORETSE_AHBo0Ii
(
CORETSE_AHBo0Ii
)
,
.CORETSE_AHBi0Ii
(
CORETSE_AHBi0Ii
)
,
.CORETSE_AHBO1Ii
(
CORETSE_AHBO1Ii
)
,
.CORETSE_AHBI1Ii
(
CORETSE_AHBI1Ii
)
,
.CORETSE_AHBl1Ii
(
CORETSE_AHBl1Ii
)
,
.CORETSE_AHBo1Ii
(
CORETSE_AHBo1Ii
)
,
.CORETSE_AHBi1Ii
(
CORETSE_AHBi1Ii
)
,
.CORETSE_AHBOoIi
(
CORETSE_AHBOoIi
)
,
.CORETSE_AHBIoIi
(
CORETSE_AHBIoIi
)
,
.CORETSE_AHBloIi
(
CORETSE_AHBloIi
)
,
.CORETSE_AHBooIi
(
CORETSE_AHBooIi
)
,
.CORETSE_AHBioIi
(
CORETSE_AHBioIi
)
,
.CORETSE_AHBOiIi
(
CORETSE_AHBOiIi
)
,
.CORETSE_AHBIiIi
(
CORETSE_AHBIiIi
)
,
.CORETSE_AHBliIi
(
CORETSE_AHBliIi
)
,
.CORETSE_AHBoiIi
(
CORETSE_AHBoiIi
)
,
.CORETSE_AHBiiIi
(
CORETSE_AHBiiIi
)
,
.CORETSE_AHBOOli
(
CORETSE_AHBOOli
)
,
.CORETSE_AHBIOli
(
CORETSE_AHBIOli
)
,
.CORETSE_AHBlOli
(
CORETSE_AHBlOli
)
,
.CORETSE_AHBoOli
(
CORETSE_AHBoOli
)
,
.CORETSE_AHBiOli
(
CORETSE_AHBiOli
)
,
.CORETSE_AHBOIli
(
CORETSE_AHBOIli
)
,
.CORETSE_AHBIIli
(
CORETSE_AHBIIli
)
,
.CORETSE_AHBlIli
(
CORETSE_AHBlIli
)
,
.CORETSE_AHBoIli
(
CORETSE_AHBoIli
)
,
.CORETSE_AHBiIli
(
CORETSE_AHBiIli
)
,
.CORETSE_AHBOlli
(
CORETSE_AHBOlli
)
,
.CORETSE_AHBIlli
(
CORETSE_AHBIlli
)
,
.CORETSE_AHBllli
(
CORETSE_AHBllli
)
,
.CORETSE_AHBolli
(
CORETSE_AHBolli
)
,
.CORETSE_AHBilli
(
CORETSE_AHBilli
)
,
.CORETSE_AHBO0li
(
CORETSE_AHBO0li
)
,
.CORETSE_AHBI0li
(
CORETSE_AHBI0li
)
,
.CORETSE_AHBl0li
(
CORETSE_AHBl0li
)
,
.CORETSE_AHBo0li
(
CORETSE_AHBo0li
)
,
.CORETSE_AHBi0li
(
CORETSE_AHBi0li
)
)
;
pemstat_eim
CORETSE_AHBo1li
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBliOi
(
CORETSE_AHBliOi
)
,
.CORETSE_AHBoiOi
(
CORETSE_AHBoiOi
)
,
.CORETSE_AHBiiOi
(
CORETSE_AHBiiOi
)
,
.CORETSE_AHBOOIi
(
CORETSE_AHBOOIi
)
,
.CORETSE_AHBooOi
(
CORETSE_AHBooOi
)
,
.CORETSE_AHBioOi
(
CORETSE_AHBioOi
)
,
.CORETSE_AHBOlIi
(
CORETSE_AHBOlIi
)
,
.CORETSE_AHBIlIi
(
CORETSE_AHBIlIi
)
,
.CORETSE_AHBllIi
(
CORETSE_AHBllIi
)
,
.CORETSE_AHBolIi
(
CORETSE_AHBolIi
)
,
.CORETSE_AHBilIi
(
CORETSE_AHBilIi
)
,
.CORETSE_AHBO0Ii
(
CORETSE_AHBO0Ii
)
,
.CORETSE_AHBI0Ii
(
CORETSE_AHBI0Ii
)
,
.CORETSE_AHBl0Ii
(
CORETSE_AHBl0Ii
)
,
.CORETSE_AHBo0Ii
(
CORETSE_AHBo0Ii
)
,
.CORETSE_AHBi0Ii
(
CORETSE_AHBi0Ii
)
,
.CORETSE_AHBO1Ii
(
CORETSE_AHBO1Ii
)
,
.CORETSE_AHBI1Ii
(
CORETSE_AHBI1Ii
)
,
.CORETSE_AHBl1Ii
(
CORETSE_AHBl1Ii
)
,
.CORETSE_AHBo1Ii
(
CORETSE_AHBo1Ii
)
,
.CORETSE_AHBi1Ii
(
CORETSE_AHBi1Ii
)
,
.CORETSE_AHBOoIi
(
CORETSE_AHBOoIi
)
,
.CORETSE_AHBIoIi
(
CORETSE_AHBIoIi
)
,
.CORETSE_AHBloIi
(
CORETSE_AHBloIi
)
,
.CORETSE_AHBooIi
(
CORETSE_AHBooIi
)
,
.CORETSE_AHBioIi
(
CORETSE_AHBioIi
)
,
.CORETSE_AHBOiIi
(
CORETSE_AHBOiIi
)
,
.CORETSE_AHBIiIi
(
CORETSE_AHBIiIi
)
,
.CORETSE_AHBliIi
(
CORETSE_AHBliIi
)
,
.CORETSE_AHBoiIi
(
CORETSE_AHBoiIi
)
,
.CORETSE_AHBiiIi
(
CORETSE_AHBiiIi
)
,
.CORETSE_AHBOOli
(
CORETSE_AHBOOli
)
,
.CORETSE_AHBIOli
(
CORETSE_AHBIOli
)
,
.CORETSE_AHBlOli
(
CORETSE_AHBlOli
)
,
.CORETSE_AHBoOli
(
CORETSE_AHBoOli
)
,
.CORETSE_AHBiOli
(
CORETSE_AHBiOli
)
,
.CORETSE_AHBOIli
(
CORETSE_AHBOIli
)
,
.CORETSE_AHBIIli
(
CORETSE_AHBIIli
)
,
.CORETSE_AHBlIli
(
CORETSE_AHBlIli
)
,
.CORETSE_AHBoIli
(
CORETSE_AHBoIli
)
,
.CORETSE_AHBiIli
(
CORETSE_AHBiIli
)
,
.CORETSE_AHBOlli
(
CORETSE_AHBOlli
)
,
.CORETSE_AHBIlli
(
CORETSE_AHBIlli
)
,
.CORETSE_AHBllli
(
CORETSE_AHBllli
)
,
.CORETSE_AHBolli
(
CORETSE_AHBolli
)
,
.CORETSE_AHBilli
(
CORETSE_AHBilli
)
,
.CORETSE_AHBO0li
(
CORETSE_AHBO0li
)
,
.CORETSE_AHBI0li
(
CORETSE_AHBI0li
)
,
.CORETSE_AHBl0li
(
CORETSE_AHBl0li
)
,
.CORETSE_AHBo0li
(
CORETSE_AHBo0li
)
,
.CORETSE_AHBi0li
(
CORETSE_AHBi0li
)
,
.CORETSE_AHBIOIi
(
CORETSE_AHBIOIi
)
,
.CORETSE_AHBlOIi
(
CORETSE_AHBlOIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBoOIi
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
)
)
;
endmodule
