// REVISION    : $Revision: 1.2 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
perex_pma
(
CORETSE_AHBIO1
,
CORETSE_AHBOO1
,
CORETSE_AHBil1
,
CORETSE_AHBlO11
,
CORETSE_AHBol1
,
CORETSE_AHBlo01
,
CORETSE_AHBlI11
,
CORETSE_AHBi010
,
CORETSE_AHBiO11
,
CORETSE_AHBOI11
)
;
input
CORETSE_AHBIO1
;
input
CORETSE_AHBOO1
;
input
[
9
:
0
]
CORETSE_AHBil1
;
input
CORETSE_AHBlO11
;
input
[
9
:
0
]
CORETSE_AHBol1
;
input
CORETSE_AHBlo01
;
input
CORETSE_AHBlI11
;
input
CORETSE_AHBi010
;
output
[
19
:
0
]
CORETSE_AHBiO11
;
output
CORETSE_AHBOI11
;
parameter
CORETSE_AHBIoII
=
1
;
reg
[
9
:
0
]
CORETSE_AHBooIOI
;
reg
[
19
:
0
]
CORETSE_AHBioIOI
;
reg
[
19
:
0
]
CORETSE_AHBOiIOI
;
wire
CORETSE_AHBIiIOI
;
wire
CORETSE_AHBliIOI
;
reg
CORETSE_AHBoiIOI
;
reg
CORETSE_AHBiiIOI
;
reg
CORETSE_AHBOOlOI
;
reg
CORETSE_AHBIOlOI
;
wire
CORETSE_AHBlOlOI
;
wire
CORETSE_AHBOI11
;
always
@
(
posedge
CORETSE_AHBIO1
or
posedge
CORETSE_AHBlI11
)
begin
if
(
CORETSE_AHBlI11
)
CORETSE_AHBooIOI
<=
#
CORETSE_AHBIoII
10
'h
0
;
else
if
(
CORETSE_AHBlo01
)
CORETSE_AHBooIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol1
;
else
CORETSE_AHBooIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBil1
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBioIOI
<=
#
CORETSE_AHBIoII
20
'h
0
;
else
if
(
CORETSE_AHBlo01
)
CORETSE_AHBioIOI
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBol1
,
CORETSE_AHBooIOI
}
;
else
CORETSE_AHBioIOI
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBil1
,
CORETSE_AHBooIOI
}
;
end
reg
[
19
:
0
]
CORETSE_AHBoOlOI
;
wire
[
9
:
0
]
CORETSE_AHBiOlOI
;
reg
[
9
:
0
]
CORETSE_AHBOIlOI
;
wire
[
19
:
0
]
CORETSE_AHBIIlOI
;
reg
[
19
:
0
]
CORETSE_AHBlIlOI
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoOlOI
<=
#
CORETSE_AHBIoII
20
'h
0
;
else
CORETSE_AHBoOlOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBioIOI
;
end
assign
CORETSE_AHBiOlOI
[
0
]
=
(
(
CORETSE_AHBoOlOI
[
6
:
0
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
6
:
0
]
==
7
'b
0000011
)
|
(
CORETSE_AHBoOlOI
[
16
:
10
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
16
:
10
]
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
1
]
=
(
(
CORETSE_AHBoOlOI
[
7
:
1
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
7
:
1
]
==
7
'b
0000011
)
|
(
CORETSE_AHBoOlOI
[
17
:
11
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
17
:
11
]
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
2
]
=
(
(
CORETSE_AHBoOlOI
[
8
:
2
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
8
:
2
]
==
7
'b
0000011
)
|
(
CORETSE_AHBoOlOI
[
18
:
12
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
18
:
12
]
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
3
]
=
(
(
CORETSE_AHBoOlOI
[
9
:
3
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
9
:
3
]
==
7
'b
0000011
)
|
(
CORETSE_AHBoOlOI
[
19
:
13
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
19
:
13
]
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
4
]
=
(
(
CORETSE_AHBoOlOI
[
10
:
4
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
10
:
4
]
==
7
'b
0000011
)
|
(
{
CORETSE_AHBioIOI
[
0
]
,
CORETSE_AHBoOlOI
[
19
:
14
]
}
==
7
'b
1111100
)
|
(
{
CORETSE_AHBioIOI
[
0
]
,
CORETSE_AHBoOlOI
[
19
:
14
]
}
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
5
]
=
(
(
CORETSE_AHBoOlOI
[
11
:
5
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
11
:
5
]
==
7
'b
0000011
)
|
(
{
CORETSE_AHBioIOI
[
1
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
15
]
}
==
7
'b
1111100
)
|
(
{
CORETSE_AHBioIOI
[
1
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
15
]
}
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
6
]
=
(
(
CORETSE_AHBoOlOI
[
12
:
6
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
12
:
6
]
==
7
'b
0000011
)
|
(
{
CORETSE_AHBioIOI
[
2
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
16
]
}
==
7
'b
1111100
)
|
(
{
CORETSE_AHBioIOI
[
2
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
16
]
}
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
7
]
=
(
(
CORETSE_AHBoOlOI
[
13
:
7
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
13
:
7
]
==
7
'b
0000011
)
|
(
{
CORETSE_AHBioIOI
[
3
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
17
]
}
==
7
'b
1111100
)
|
(
{
CORETSE_AHBioIOI
[
3
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
17
]
}
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
8
]
=
(
(
CORETSE_AHBoOlOI
[
14
:
8
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
14
:
8
]
==
7
'b
0000011
)
|
(
{
CORETSE_AHBioIOI
[
4
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
18
]
}
==
7
'b
1111100
)
|
(
{
CORETSE_AHBioIOI
[
4
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
18
]
}
==
7
'b
0000011
)
)
;
assign
CORETSE_AHBiOlOI
[
9
]
=
(
(
CORETSE_AHBoOlOI
[
15
:
9
]
==
7
'b
1111100
)
|
(
CORETSE_AHBoOlOI
[
15
:
9
]
==
7
'b
0000011
)
|
(
{
CORETSE_AHBioIOI
[
5
:
0
]
,
CORETSE_AHBoOlOI
[
19
]
}
==
7
'b
1111100
)
|
(
{
CORETSE_AHBioIOI
[
5
:
0
]
,
CORETSE_AHBoOlOI
[
19
]
}
==
7
'b
0000011
)
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOIlOI
<=
#
CORETSE_AHBIoII
10
'h
001
;
else
if
(
|
CORETSE_AHBiOlOI
)
CORETSE_AHBOIlOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOlOI
;
end
assign
CORETSE_AHBIIlOI
=
{
20
{
CORETSE_AHBOIlOI
==
10
'h
001
}
}
&
CORETSE_AHBoOlOI
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
1
]
==
9
'h
001
}
}
&
{
CORETSE_AHBioIOI
[
0
]
,
CORETSE_AHBoOlOI
[
19
:
1
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
2
]
==
8
'h
01
}
}
&
{
CORETSE_AHBioIOI
[
1
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
2
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
3
]
==
7
'h
01
}
}
&
{
CORETSE_AHBioIOI
[
2
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
3
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
4
]
==
6
'h
01
}
}
&
{
CORETSE_AHBioIOI
[
3
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
4
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
5
]
==
5
'h
01
}
}
&
{
CORETSE_AHBioIOI
[
4
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
5
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
6
]
==
4
'h
1
}
}
&
{
CORETSE_AHBioIOI
[
5
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
6
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
7
]
==
3
'h
1
}
}
&
{
CORETSE_AHBioIOI
[
6
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
7
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
:
8
]
==
2
'h
1
}
}
&
{
CORETSE_AHBioIOI
[
7
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
8
]
}
|
{
20
{
CORETSE_AHBOIlOI
[
9
]
==
1
'b
1
}
}
&
{
CORETSE_AHBioIOI
[
8
:
0
]
,
CORETSE_AHBoOlOI
[
19
:
9
]
}
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlIlOI
<=
#
CORETSE_AHBIoII
20
'h
0
;
else
CORETSE_AHBlIlOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIlOI
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOiIOI
<=
#
CORETSE_AHBIoII
20
'h
0
;
else
CORETSE_AHBOiIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIlOI
;
end
assign
CORETSE_AHBIiIOI
=
CORETSE_AHBlIlOI
[
9
:
0
]
==
10
'b
01_0111_1100
|
CORETSE_AHBlIlOI
[
9
:
0
]
==
10
'b
10_1000_0011
|
CORETSE_AHBlIlOI
[
9
:
0
]
==
10
'b
10_0111_1100
|
CORETSE_AHBlIlOI
[
9
:
0
]
==
10
'b
01_1000_0011
;
assign
CORETSE_AHBliIOI
=
CORETSE_AHBlIlOI
[
19
:
10
]
==
10
'b
01_0111_1100
|
CORETSE_AHBlIlOI
[
19
:
10
]
==
10
'b
10_1000_0011
|
CORETSE_AHBlIlOI
[
19
:
10
]
==
10
'b
10_0111_1100
|
CORETSE_AHBlIlOI
[
19
:
10
]
==
10
'b
01_1000_0011
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoiIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoiIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIiIOI
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiiIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiiIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBliIOI
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOOlOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOOlOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiIOI
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIOlOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBlO11
)
CORETSE_AHBIOlOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBliIOI
&
~
CORETSE_AHBIiIOI
)
CORETSE_AHBIOlOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBIiIOI
&
~
CORETSE_AHBliIOI
)
CORETSE_AHBIOlOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
assign
CORETSE_AHBiO11
=
{
20
{
CORETSE_AHBIOlOI
}
}
&
CORETSE_AHBOiIOI
|
{
20
{
~
CORETSE_AHBIOlOI
}
}
&
{
CORETSE_AHBlIlOI
[
9
:
0
]
,
CORETSE_AHBOiIOI
[
19
:
10
]
}
;
assign
CORETSE_AHBlOlOI
=
(
CORETSE_AHBIOlOI
&
(
(
CORETSE_AHBiiIOI
&
CORETSE_AHBoiIOI
)
|
(
CORETSE_AHBOOlOI
&
CORETSE_AHBoiIOI
)
)
)
|
(
~
CORETSE_AHBIOlOI
&
(
(
CORETSE_AHBIiIOI
&
CORETSE_AHBiiIOI
)
|
(
CORETSE_AHBiiIOI
&
CORETSE_AHBoiIOI
)
)
)
;
assign
CORETSE_AHBOI11
=
1
'b
0
;
endmodule
