// REVISION    : $Revision: 1.6 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxrfif_fab
#
(
parameter
RABITS
=
12
,
parameter
CORETSE_AHBIo1
=
32
,
parameter
CORETSE_AHBlo1
=
$clog2
(
CORETSE_AHBIo1
/
8
)
)
(
CORETSE_AHBOlo
,
CORETSE_AHBI0II
,
CORETSE_AHBIOII
,
CORETSE_AHBIlo
,
CORETSE_AHBi0i
,
CORETSE_AHBIii
,
CORETSE_AHBlii
,
CORETSE_AHBoii
,
CORETSE_AHBllII
,
CORETSE_AHBolII
,
CORETSE_AHBOIOI
,
CORETSE_AHBo0i
,
CORETSE_AHBioo
,
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBoio
,
CORETSE_AHBooi
,
CORETSE_AHBioi
,
CORETSE_AHBOii
,
CORETSE_AHBO0OI
,
CORETSE_AHBI0OI
)
;
input
CORETSE_AHBOlo
;
input
CORETSE_AHBI0II
;
input
CORETSE_AHBIOII
;
input
CORETSE_AHBIlo
;
input
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBi0i
;
input
[
RABITS
:
0
]
CORETSE_AHBIii
;
input
CORETSE_AHBlii
;
input
CORETSE_AHBoii
;
input
[
RABITS
+
1
:
0
]
CORETSE_AHBllII
;
input
CORETSE_AHBolII
;
output
CORETSE_AHBOIOI
;
output
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBo0i
;
output
[
(
CORETSE_AHBIo1
-
1
)
:
0
]
CORETSE_AHBioo
;
output
CORETSE_AHBOio
;
output
CORETSE_AHBIio
;
output
[
1
:
0
]
CORETSE_AHBlio
;
output
CORETSE_AHBoio
;
output
CORETSE_AHBooi
;
output
[
RABITS
:
0
]
CORETSE_AHBioi
;
output
CORETSE_AHBOii
;
output
CORETSE_AHBO0OI
;
output
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBI0OI
;
parameter
CORETSE_AHBol0I
=
{
(
RABITS
+
1
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBIoII
=
1
;
wire
CORETSE_AHBil0I
;
reg
CORETSE_AHBO00I
;
reg
[
RABITS
:
0
]
CORETSE_AHBI00I
;
wire
[
RABITS
:
0
]
CORETSE_AHBl00I
;
wire
[
RABITS
:
0
]
CORETSE_AHBo00I
;
reg
[
RABITS
:
0
]
CORETSE_AHBi00I
;
reg
CORETSE_AHBOIOI
;
reg
CORETSE_AHBO10I
;
reg
CORETSE_AHBooi
;
reg
CORETSE_AHBOii
;
reg
[
RABITS
:
0
]
CORETSE_AHBioi
;
reg
CORETSE_AHBI10I
,
CORETSE_AHBl10I
;
reg
CORETSE_AHBo10I
,
CORETSE_AHBi10I
;
reg
CORETSE_AHBOo0I
,
CORETSE_AHBIo0I
;
reg
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBlo0I
;
reg
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBoo0I
;
reg
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBio0I
;
reg
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBOi0I
;
reg
[
3
:
0
]
CORETSE_AHBIi0I
;
wire
CORETSE_AHBoio
;
reg
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBI0OI
;
reg
CORETSE_AHBO0OI
;
reg
CORETSE_AHBli0I
;
reg
CORETSE_AHBoi0I
;
reg
CORETSE_AHBii0I
;
wire
CORETSE_AHBOO1I
;
wire
CORETSE_AHBIO1I
;
//      generate logic as part of synthesis results.
wire
[
(
RABITS
-
1
)
:
0
]
#
1000
CORETSE_AHBo0i
=
(
{
RABITS
{
~
(
~
CORETSE_AHBllII
[
RABITS
+
1
]
&
CORETSE_AHBOO1I
)
}
}
&
(
CORETSE_AHBl00I
[
(
RABITS
-
1
)
:
0
]
-
'd
1
)
)
|
(
{
RABITS
{
(
~
CORETSE_AHBllII
[
RABITS
+
1
]
&
CORETSE_AHBOO1I
)
}
}
&
(
CORETSE_AHBllII
[
(
RABITS
-
1
)
:
0
]
)
)
;
assign
CORETSE_AHBo00I
=
CORETSE_AHBi00I
+
1
'b
1
;
assign
CORETSE_AHBil0I
=
(
(
CORETSE_AHBI00I
[
RABITS
:
0
]
!=
CORETSE_AHBi00I
[
RABITS
:
0
]
)
&
CORETSE_AHBOIOI
&
~
CORETSE_AHBIi0I
[
1
]
)
;
assign
CORETSE_AHBl00I
=
CORETSE_AHBil0I
?
CORETSE_AHBo00I
:
CORETSE_AHBi00I
;
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBi00I
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
CORETSE_AHBi00I
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBO00I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO00I
<=
#
CORETSE_AHBIoII
CORETSE_AHBil0I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
begin
CORETSE_AHBlo0I
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
4
)
{
1
'b
0
}
}
;
CORETSE_AHBoo0I
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
4
)
{
1
'b
0
}
}
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
4
)
{
1
'b
0
}
}
;
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
4
)
{
1
'b
0
}
}
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
0
;
end
else
begin
case
(
{
CORETSE_AHBIlo
,
CORETSE_AHBO00I
,
CORETSE_AHBIi0I
}
)
6
'b
010000
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
8
;
end
6
'b
011000
:
begin
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
C
;
end
6
'b
011100
:
begin
CORETSE_AHBoo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
E
;
end
6
'b
011110
:
begin
CORETSE_AHBlo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
F
;
end
6
'b
101000
:
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
0
;
6
'b
101100
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
8
;
end
6
'b
101110
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0I
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
C
;
end
6
'b
101111
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0I
;
CORETSE_AHBoo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo0I
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
E
;
end
6
'b
110000
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
4
'h
8
;
end
6
'b
111000
:
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
6
'b
111100
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
end
6
'b
111110
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0I
;
CORETSE_AHBoo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
end
6
'b
111111
:
begin
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0I
;
CORETSE_AHBoo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo0I
;
CORETSE_AHBlo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0i
;
end
default
:
begin
CORETSE_AHBlo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo0I
;
CORETSE_AHBoo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0I
;
CORETSE_AHBio0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBio0I
;
CORETSE_AHBOi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi0I
;
CORETSE_AHBIi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi0I
;
end
endcase
end
end
assign
{
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBioo
}
=
CORETSE_AHBOi0I
;
assign
CORETSE_AHBoio
=
CORETSE_AHBIi0I
[
3
]
;
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBO10I
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
if
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
&
CORETSE_AHBOio
)
CORETSE_AHBO10I
<=
#
CORETSE_AHBIoII
1
'h
1
;
else
if
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
&
CORETSE_AHBIio
)
CORETSE_AHBO10I
<=
#
CORETSE_AHBIoII
1
'h
0
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBOIOI
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
if
(
CORETSE_AHBOo0I
)
CORETSE_AHBOIOI
<=
#
CORETSE_AHBIoII
1
'h
1
;
else
if
(
~
CORETSE_AHBO10I
&
(
CORETSE_AHBI00I
[
RABITS
:
0
]
!=
CORETSE_AHBi00I
[
RABITS
:
0
]
)
)
CORETSE_AHBOIOI
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOIOI
<=
#
CORETSE_AHBIoII
1
'h
0
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBOii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo10I
)
CORETSE_AHBOii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOii
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBioi
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
~
CORETSE_AHBOii
&
~
CORETSE_AHBo10I
)
CORETSE_AHBioi
<=
#
CORETSE_AHBIoII
CORETSE_AHBi00I
[
RABITS
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBooi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
~
CORETSE_AHBI10I
)
CORETSE_AHBooi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBI10I
)
CORETSE_AHBooi
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBI00I
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBI10I
&
~
CORETSE_AHBooi
)
CORETSE_AHBI00I
<=
#
CORETSE_AHBIoII
CORETSE_AHBIii
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBi10I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi10I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoii
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBo10I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo10I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi10I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBl10I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl10I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlii
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBI10I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI10I
<=
#
CORETSE_AHBIoII
CORETSE_AHBl10I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBli0I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBli0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBolII
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBoi0I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoi0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBli0I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBii0I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBii0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoi0I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBO0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBii0I
;
end
assign
CORETSE_AHBOO1I
=
CORETSE_AHBoi0I
&
~
CORETSE_AHBii0I
;
assign
CORETSE_AHBIO1I
=
CORETSE_AHBii0I
&
~
CORETSE_AHBO0OI
;
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBI0OI
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
{
1
'b
0
}
}
;
else
if
(
~
CORETSE_AHBllII
[
RABITS
+
1
]
&
CORETSE_AHBIO1I
)
CORETSE_AHBI0OI
<=
#
CORETSE_AHBIoII
{
{
(
CORETSE_AHBlo1
+
2
)
{
1
'b
0
}
}
,
CORETSE_AHBi0i
}
;
else
if
(
CORETSE_AHBllII
[
RABITS
+
1
]
&
CORETSE_AHBOO1I
)
CORETSE_AHBI0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00I
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBIo0I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOII
;
end
always
@
(
posedge
CORETSE_AHBOlo
or
posedge
CORETSE_AHBI0II
)
begin
if
(
CORETSE_AHBI0II
)
CORETSE_AHBOo0I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOo0I
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo0I
;
end
endmodule
