// REVISION    : $Revision: 1.6 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
pehst
(
CORETSE_AHBio1
,
CORETSE_AHBOi1
,
CORETSE_AHBIi1
,
CORETSE_AHBli1
,
CORETSE_AHBoi1
,
CORETSE_AHBii1
,
CORETSE_AHBOi11
,
CORETSE_AHBOIi1
,
CORETSE_AHBiOi1
,
CORETSE_AHBIIi1
,
CORETSE_AHBlIi1
,
CORETSE_AHBiIi
,
CORETSE_AHBIOi1
,
CORETSE_AHBlOi1
,
CORETSE_AHBoOi1
,
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
,
CORETSE_AHBI000
,
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
,
CORETSE_AHBO1i
,
CORETSE_AHBI1i
,
CORETSE_AHBoIi1
,
CORETSE_AHBiIi1
,
CORETSE_AHBll00
,
CORETSE_AHBOoOo
,
CORETSE_AHBi111
,
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
,
CORETSE_AHBio01
,
CORETSE_AHBi0i1
,
CORETSE_AHBO1i1
,
CORETSE_AHBI1i1
,
CORETSE_AHBIii1
,
CORETSE_AHBOii1
,
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
,
CORETSE_AHBi1i1
,
CORETSE_AHBOoi1
,
CORETSE_AHBoii1
,
CORETSE_AHBiii1
,
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
,
CORETSE_AHBooi1
,
CORETSE_AHBioi1
,
CORETSE_AHBoiOo
,
CORETSE_AHBoo01
,
CORETSE_AHBOli1
,
CORETSE_AHBIli1
,
CORETSE_AHBlli1
,
CORETSE_AHBlii1
,
CORETSE_AHBOOOo
,
CORETSE_AHBIOOo
,
CORETSE_AHBiii0
,
CORETSE_AHBlOOo
,
CORETSE_AHBoOOo
,
CORETSE_AHBiOOo
,
CORETSE_AHBOIOo
,
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
,
CORETSE_AHBIIOo
,
CORETSE_AHBlIOo
,
CORETSE_AHBoIOo
,
CORETSE_AHBiIOo
,
CORETSE_AHBOlOo
,
CORETSE_AHBIlOo
,
CORETSE_AHBii01
,
CORETSE_AHBllOo
,
CORETSE_AHBolOo
,
CORETSE_AHBilOo
,
CORETSE_AHBO0Oo
,
CORETSE_AHBI0Oo
,
CORETSE_AHBiiOo
,
CORETSE_AHBl0Oo
,
CORETSE_AHBOOIo
,
CORETSE_AHBIOIo
)
;
input
CORETSE_AHBio1
,
CORETSE_AHBOi1
,
CORETSE_AHBIi1
,
CORETSE_AHBli1
;
input
[
7
:
0
]
CORETSE_AHBoi1
;
input
[
31
:
0
]
CORETSE_AHBii1
;
input
[
4
:
0
]
CORETSE_AHBOi11
;
input
[
15
:
0
]
CORETSE_AHBOIi1
;
input
CORETSE_AHBiOi1
,
CORETSE_AHBIIi1
,
CORETSE_AHBlIi1
;
input
CORETSE_AHBiIi
;
input
CORETSE_AHBIOi1
,
CORETSE_AHBlOi1
;
input
CORETSE_AHBoOi1
;
input
CORETSE_AHBI000
;
output
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
;
output
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
;
output
[
31
:
0
]
CORETSE_AHBO1i
;
output
CORETSE_AHBI1i
;
output
CORETSE_AHBoIi1
,
CORETSE_AHBiIi1
;
output
[
47
:
0
]
CORETSE_AHBll00
;
output
[
15
:
0
]
CORETSE_AHBOoOo
;
output
[
15
:
0
]
CORETSE_AHBi111
;
output
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
;
output
CORETSE_AHBio01
,
CORETSE_AHBi0i1
,
CORETSE_AHBO1i1
;
output
[
6
:
0
]
CORETSE_AHBI1i1
;
output
[
7
:
0
]
CORETSE_AHBIii1
;
output
[
15
:
0
]
CORETSE_AHBOii1
;
output
[
6
:
0
]
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
;
output
[
3
:
0
]
CORETSE_AHBoii1
;
output
CORETSE_AHBiii1
;
output
[
9
:
0
]
CORETSE_AHBi1i1
;
output
[
3
:
0
]
CORETSE_AHBOoi1
;
output
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
;
output
CORETSE_AHBOli1
,
CORETSE_AHBIli1
,
CORETSE_AHBlli1
;
output
CORETSE_AHBooi1
,
CORETSE_AHBioi1
;
output
[
1
:
0
]
CORETSE_AHBoo01
;
output
CORETSE_AHBoiOo
;
output
[
3
:
0
]
CORETSE_AHBlii1
;
output
CORETSE_AHBOOOo
,
CORETSE_AHBIOOo
;
output
CORETSE_AHBiii0
,
CORETSE_AHBlOOo
;
output
[
2
:
0
]
CORETSE_AHBoOOo
;
output
CORETSE_AHBiOOo
,
CORETSE_AHBOIOo
;
output
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
;
output
[
4
:
0
]
CORETSE_AHBIIOo
,
CORETSE_AHBlIOo
;
output
CORETSE_AHBoIOo
;
output
[
15
:
0
]
CORETSE_AHBiIOo
;
output
CORETSE_AHBOlOo
,
CORETSE_AHBIlOo
;
output
CORETSE_AHBii01
;
output
CORETSE_AHBllOo
,
CORETSE_AHBolOo
,
CORETSE_AHBilOo
,
CORETSE_AHBO0Oo
;
output
CORETSE_AHBI0Oo
;
output
CORETSE_AHBiiOo
,
CORETSE_AHBl0Oo
;
output
CORETSE_AHBOOIo
,
CORETSE_AHBIOIo
;
wire
[
31
:
0
]
CORETSE_AHBO1i
;
wire
CORETSE_AHBI1i
;
reg
CORETSE_AHBoIi1
,
CORETSE_AHBiIi1
;
reg
[
47
:
0
]
CORETSE_AHBll00
;
reg
[
15
:
0
]
CORETSE_AHBOoOo
;
reg
[
15
:
0
]
CORETSE_AHBi111
;
reg
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
;
reg
CORETSE_AHBio01
,
CORETSE_AHBi0i1
,
CORETSE_AHBO1i1
;
reg
[
6
:
0
]
CORETSE_AHBI1i1
;
reg
[
15
:
0
]
CORETSE_AHBOii1
;
reg
[
7
:
0
]
CORETSE_AHBIii1
;
reg
[
6
:
0
]
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
;
reg
[
3
:
0
]
CORETSE_AHBoii1
;
reg
CORETSE_AHBiii1
;
reg
[
9
:
0
]
CORETSE_AHBi1i1
;
reg
[
3
:
0
]
CORETSE_AHBOoi1
;
reg
CORETSE_AHBOli1
,
CORETSE_AHBIli1
,
CORETSE_AHBlli1
;
reg
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
;
wire
CORETSE_AHBooi1
;
reg
CORETSE_AHBioi1
;
reg
[
1
:
0
]
CORETSE_AHBoo01
;
reg
CORETSE_AHBoiOo
;
reg
[
3
:
0
]
CORETSE_AHBlii1
;
reg
CORETSE_AHBOOOo
,
CORETSE_AHBIOOo
;
reg
CORETSE_AHBiii0
,
CORETSE_AHBlOOo
;
reg
[
2
:
0
]
CORETSE_AHBoOOo
;
reg
CORETSE_AHBiOOo
,
CORETSE_AHBOIOo
;
reg
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
;
reg
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
;
reg
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
;
reg
[
4
:
0
]
CORETSE_AHBIIOo
,
CORETSE_AHBlIOo
;
wire
CORETSE_AHBoIOo
;
reg
[
15
:
0
]
CORETSE_AHBiIOo
;
reg
CORETSE_AHBOlOo
,
CORETSE_AHBIlOo
;
reg
CORETSE_AHBii01
;
reg
CORETSE_AHBllOo
,
CORETSE_AHBolOo
,
CORETSE_AHBilOo
,
CORETSE_AHBO0Oo
;
reg
CORETSE_AHBI0Oo
;
reg
CORETSE_AHBiiOo
,
CORETSE_AHBl0Oo
;
reg
CORETSE_AHBOOIo
,
CORETSE_AHBIOIo
;
parameter
CORETSE_AHBIoII
=
1
;
wire
CORETSE_AHBl11o
,
CORETSE_AHBo11o
;
wire
CORETSE_AHBi11o
,
CORETSE_AHBOo1o
;
reg
CORETSE_AHBIo1o
;
wire
CORETSE_AHBlo1o
,
CORETSE_AHBoo1o
;
wire
CORETSE_AHBio1o
,
CORETSE_AHBOi1o
;
wire
CORETSE_AHBIi1o
,
CORETSE_AHBli1o
;
wire
CORETSE_AHBoi1o
,
CORETSE_AHBii1o
;
wire
CORETSE_AHBOOoo
,
CORETSE_AHBIOoo
;
wire
CORETSE_AHBlOoo
,
CORETSE_AHBoOoo
;
wire
CORETSE_AHBiOoo
;
wire
CORETSE_AHBOIoo
,
CORETSE_AHBIIoo
;
wire
CORETSE_AHBlIoo
,
CORETSE_AHBoIoo
;
wire
CORETSE_AHBiIoo
,
CORETSE_AHBOloo
;
wire
CORETSE_AHBIloo
,
CORETSE_AHBlloo
;
wire
CORETSE_AHBoloo
;
wire
CORETSE_AHBiloo
;
wire
CORETSE_AHBO0oo
;
reg
CORETSE_AHBI0oo
;
reg
CORETSE_AHBl0oo
,
CORETSE_AHBo0oo
,
CORETSE_AHBi0oo
;
wire
CORETSE_AHBO1oo
;
reg
CORETSE_AHBI1oo
,
CORETSE_AHBl1oo
,
CORETSE_AHBo1oo
;
wire
CORETSE_AHBi1oo
,
CORETSE_AHBOooo
;
wire
CORETSE_AHBIooo
,
CORETSE_AHBlooo
;
assign
CORETSE_AHBl11o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
00
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBo11o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
00
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBi11o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
01
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOo1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
01
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBlo1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
02
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoo1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
02
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBio1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
03
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOi1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
03
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBIi1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
04
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBli1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
04
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoi1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
05
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBii1o
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
05
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOOoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
06
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBIOoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
06
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOIoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
07
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBIIoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
07
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBlIoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
08
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoIoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
08
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBiIoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
09
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOloo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
09
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBIloo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0a
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBlloo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0a
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoIOo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0b
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoloo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0b
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBiloo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0c
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBO0oo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0d
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBlOoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0e
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoOoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0e
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBiOoo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
0f
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBi1oo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
10
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOooo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
10
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBIooo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
11
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBlooo
=
CORETSE_AHBoi1
[
7
:
0
]
==
8
'h
11
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBii01
,
CORETSE_AHBlOOo
,
CORETSE_AHBO0Oo
,
CORETSE_AHBilOo
,
CORETSE_AHBolOo
,
CORETSE_AHBllOo
,
CORETSE_AHBiii0
,
CORETSE_AHBiIi1
,
CORETSE_AHBoIi1
,
CORETSE_AHBOOOo
,
CORETSE_AHBIOOo
}
<=
#
CORETSE_AHBIoII
{
2
'b
10
,
4
'b
0000
,
1
'b
0
,
2
'b
00
,
2
'b
00
}
;
else
if
(
CORETSE_AHBl11o
)
{
CORETSE_AHBii01
,
CORETSE_AHBlOOo
,
CORETSE_AHBO0Oo
,
CORETSE_AHBilOo
,
CORETSE_AHBolOo
,
CORETSE_AHBllOo
,
CORETSE_AHBiii0
,
CORETSE_AHBiIi1
,
CORETSE_AHBoIi1
,
CORETSE_AHBOOOo
,
CORETSE_AHBIOOo
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
:
30
]
,
CORETSE_AHBii1
[
19
:
16
]
,
CORETSE_AHBii1
[
8
]
,
CORETSE_AHBii1
[
5
:
4
]
,
CORETSE_AHBii1
[
2
]
,
CORETSE_AHBii1
[
0
]
}
;
end
assign
CORETSE_AHBooi1
=
CORETSE_AHBiIi
|
CORETSE_AHBIo1o
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBlii1
,
CORETSE_AHBoo01
,
CORETSE_AHBO1i1
,
CORETSE_AHBi0i1
,
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
,
CORETSE_AHBio01
}
<=
#
CORETSE_AHBIoII
{
4
'b
0111
,
2
'b
10
,
2
'b
00
,
3
'b
000
}
;
else
if
(
CORETSE_AHBi11o
)
{
CORETSE_AHBlii1
,
CORETSE_AHBoo01
,
CORETSE_AHBO1i1
,
CORETSE_AHBi0i1
,
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
,
CORETSE_AHBio01
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
15
:
12
]
,
CORETSE_AHBii1
[
9
:
8
]
,
CORETSE_AHBii1
[
5
:
4
]
,
CORETSE_AHBii1
[
2
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
,
CORETSE_AHBIii1
,
CORETSE_AHBI1i1
}
<=
#
CORETSE_AHBIoII
{
7
'h
40
,
7
'h
60
,
8
'h
50
,
7
'h
60
}
;
else
if
(
CORETSE_AHBlo1o
)
{
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
,
CORETSE_AHBIii1
,
CORETSE_AHBI1i1
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
30
:
24
]
,
CORETSE_AHBii1
[
22
:
16
]
,
CORETSE_AHBii1
[
15
:
8
]
,
CORETSE_AHBii1
[
6
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBoii1
,
CORETSE_AHBiii1
,
CORETSE_AHBioi1
,
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
,
CORETSE_AHBOoi1
,
CORETSE_AHBi1i1
}
<=
#
CORETSE_AHBIoII
{
4
'h
a
,
4
'b
0001
,
4
'h
f
,
10
'h
37
}
;
else
if
(
CORETSE_AHBio1o
)
{
CORETSE_AHBoii1
,
CORETSE_AHBiii1
,
CORETSE_AHBioi1
,
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
,
CORETSE_AHBOoi1
,
CORETSE_AHBi1i1
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
23
:
20
]
,
CORETSE_AHBii1
[
19
:
16
]
,
CORETSE_AHBii1
[
15
:
12
]
,
CORETSE_AHBii1
[
9
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBI1oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI1oo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi1o
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBl1oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1oo
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1oo
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBo1oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo1oo
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1oo
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBOii1
<=
#
CORETSE_AHBIoII
16
'h
07D0
;
else
if
(
CORETSE_AHBIi1o
)
CORETSE_AHBOii1
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBOoOo
<=
#
CORETSE_AHBIoII
16
'h
0000
;
else
if
(
CORETSE_AHBoi1o
)
CORETSE_AHBOoOo
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBi111
<=
#
CORETSE_AHBIoII
16
'h
FFFF
;
else
if
(
CORETSE_AHBOOoo
)
CORETSE_AHBi111
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBlli1
,
CORETSE_AHBIo1o
,
CORETSE_AHBOli1
,
CORETSE_AHBIli1
}
<=
#
CORETSE_AHBIoII
4
'h
0
;
else
if
(
CORETSE_AHBOIoo
)
{
CORETSE_AHBlli1
,
CORETSE_AHBIo1o
,
CORETSE_AHBOli1
,
CORETSE_AHBIli1
}
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
3
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBI0Oo
,
CORETSE_AHBOIOo
,
CORETSE_AHBiOOo
,
CORETSE_AHBoOOo
}
<=
#
CORETSE_AHBIoII
6
'h
00
;
else
if
(
CORETSE_AHBlIoo
)
{
CORETSE_AHBI0Oo
,
CORETSE_AHBOIOo
,
CORETSE_AHBiOOo
,
CORETSE_AHBoOOo
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
]
,
CORETSE_AHBii1
[
5
:
4
]
,
CORETSE_AHBii1
[
2
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBIlOo
,
CORETSE_AHBOlOo
}
<=
#
CORETSE_AHBIoII
2
'h
0
;
else
if
(
CORETSE_AHBiIoo
)
{
CORETSE_AHBIlOo
,
CORETSE_AHBOlOo
}
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
1
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBIIOo
,
CORETSE_AHBlIOo
}
<=
#
CORETSE_AHBIoII
{
5
'h
0
,
5
'h
0
}
;
else
if
(
CORETSE_AHBIloo
)
{
CORETSE_AHBIIOo
,
CORETSE_AHBlIOo
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
12
:
8
]
,
CORETSE_AHBii1
[
4
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBiIOo
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBoIOo
)
CORETSE_AHBiIOo
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBl0Oo
,
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
,
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
,
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
}
<=
#
CORETSE_AHBIoII
13
'h
0
;
else
if
(
CORETSE_AHBlOoo
)
{
CORETSE_AHBl0Oo
,
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
,
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
,
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
]
,
CORETSE_AHBii1
[
27
:
25
]
,
CORETSE_AHBii1
[
7
:
4
]
,
CORETSE_AHBii1
[
3
:
2
]
}
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBI0oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBIIi1
)
CORETSE_AHBI0oo
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBO1oo
)
CORETSE_AHBI0oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBl0oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl0oo
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOoo
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBo0oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo0oo
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0oo
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBi0oo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi0oo
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0oo
;
end
assign
CORETSE_AHBO1oo
=
~
CORETSE_AHBo0oo
&
CORETSE_AHBi0oo
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBll00
[
7
:
0
]
,
CORETSE_AHBll00
[
15
:
8
]
,
CORETSE_AHBll00
[
23
:
16
]
,
CORETSE_AHBll00
[
31
:
24
]
}
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
if
(
CORETSE_AHBi1oo
)
{
CORETSE_AHBll00
[
7
:
0
]
,
CORETSE_AHBll00
[
15
:
8
]
,
CORETSE_AHBll00
[
23
:
16
]
,
CORETSE_AHBll00
[
31
:
24
]
}
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
31
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBll00
[
39
:
32
]
,
CORETSE_AHBll00
[
47
:
40
]
}
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBIooo
)
{
CORETSE_AHBll00
[
39
:
32
]
,
CORETSE_AHBll00
[
47
:
40
]
}
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
31
:
16
]
;
end
assign
CORETSE_AHBI1i
=
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBO1i
[
31
:
0
]
=
{
32
{
CORETSE_AHBlooo
}
}
&
{
CORETSE_AHBll00
[
39
:
32
]
,
CORETSE_AHBll00
[
47
:
40
]
,
16
'h
0
}
|
{
32
{
CORETSE_AHBOooo
}
}
&
{
CORETSE_AHBll00
[
7
:
0
]
,
CORETSE_AHBll00
[
15
:
8
]
,
CORETSE_AHBll00
[
23
:
16
]
,
CORETSE_AHBll00
[
31
:
24
]
}
|
{
32
{
CORETSE_AHBiOoo
}
}
&
{
21
'h
0
,
CORETSE_AHBI000
,
CORETSE_AHBoOi1
,
5
'b
0
,
CORETSE_AHBI0oo
,
3
'b
0
}
|
{
32
{
CORETSE_AHBoOoo
}
}
&
{
CORETSE_AHBl0Oo
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
,
1
'b
0
,
16
'b
0
,
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
,
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
,
2
'b
0
}
|
{
32
{
CORETSE_AHBO0oo
}
}
&
{
16
'h
0
,
13
'h
0
,
CORETSE_AHBlIi1
,
CORETSE_AHBIlOo
,
CORETSE_AHBiOi1
}
|
{
32
{
CORETSE_AHBiloo
}
}
&
{
16
'h
0
,
CORETSE_AHBOIi1
[
15
:
0
]
}
|
{
32
{
CORETSE_AHBoloo
}
}
&
{
16
'h
0
,
CORETSE_AHBiIOo
[
15
:
0
]
}
|
{
32
{
CORETSE_AHBlloo
}
}
&
{
16
'h
0
,
3
'h
0
,
CORETSE_AHBIIOo
[
4
:
0
]
,
3
'h
0
,
CORETSE_AHBlIOo
[
4
:
0
]
}
|
{
32
{
CORETSE_AHBOloo
}
}
&
{
28
'h
0
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBIlOo
,
CORETSE_AHBOlOo
}
|
{
32
{
CORETSE_AHBoIoo
}
}
&
{
CORETSE_AHBI0Oo
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
20
'h
0
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBOIOo
,
CORETSE_AHBiOOo
,
1
'b
0
,
CORETSE_AHBoOOo
[
2
:
0
]
}
|
{
32
{
CORETSE_AHBIIoo
}
}
&
{
16
'h
0
,
12
'h
0
,
CORETSE_AHBlli1
,
CORETSE_AHBIo1o
,
CORETSE_AHBOli1
,
CORETSE_AHBIli1
}
|
{
32
{
CORETSE_AHBli1o
}
}
&
{
16
'h
0
,
CORETSE_AHBOii1
[
15
:
0
]
}
|
{
32
{
CORETSE_AHBii1o
}
}
&
{
16
'h
0
,
CORETSE_AHBOoOo
[
15
:
0
]
}
|
{
32
{
CORETSE_AHBIOoo
}
}
&
{
16
'h
0
,
CORETSE_AHBi111
[
15
:
0
]
}
|
{
32
{
CORETSE_AHBOi1o
}
}
&
{
8
'h
0
,
CORETSE_AHBoii1
[
3
:
0
]
,
CORETSE_AHBiii1
,
CORETSE_AHBioi1
,
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
,
CORETSE_AHBOoi1
[
3
:
0
]
,
2
'h
0
,
CORETSE_AHBi1i1
[
9
:
0
]
}
|
{
32
{
CORETSE_AHBoo1o
}
}
&
{
1
'b
0
,
CORETSE_AHBl1i1
[
6
:
0
]
,
1
'b
0
,
CORETSE_AHBo1i1
[
6
:
0
]
,
CORETSE_AHBIii1
[
7
:
0
]
,
1
'b
0
,
CORETSE_AHBI1i1
[
6
:
0
]
}
|
{
32
{
CORETSE_AHBOo1o
}
}
&
{
16
'h
0
,
CORETSE_AHBlii1
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBoo01
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBO1i1
,
CORETSE_AHBi0i1
,
1
'b
0
,
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
,
CORETSE_AHBio01
}
|
{
32
{
CORETSE_AHBo11o
}
}
&
{
CORETSE_AHBii01
,
CORETSE_AHBlOOo
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBO0Oo
,
CORETSE_AHBilOo
,
CORETSE_AHBolOo
,
CORETSE_AHBllOo
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBiii0
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBiIi1
,
CORETSE_AHBoIi1
,
CORETSE_AHBIOi1
,
CORETSE_AHBOOOo
,
CORETSE_AHBlOi1
,
CORETSE_AHBIOOo
}
;
endmodule
