// REVISION    : $Revision: 1.3 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxtfif_wtm
#
(
parameter
RABITS
=
12
)
(
CORETSE_AHBoi0
,
CORETSE_AHBllo
,
CORETSE_AHBo0II
,
CORETSE_AHBoOII
,
CORETSE_AHBl0OI
,
CORETSE_AHBo0OI
,
CORETSE_AHBi0OI
,
CORETSE_AHBO1OI
,
CORETSE_AHBI1OI
,
CORETSE_AHBIoo
,
CORETSE_AHBiii
,
CORETSE_AHBIOOI
,
CORETSE_AHBOOOI
,
CORETSE_AHBlIOI
,
CORETSE_AHBlIi
,
CORETSE_AHBoIi
,
CORETSE_AHBiIi
,
CORETSE_AHBlOOI
)
;
input
CORETSE_AHBoi0
;
input
CORETSE_AHBllo
;
input
CORETSE_AHBo0II
;
input
CORETSE_AHBoOII
;
input
[
15
:
0
]
CORETSE_AHBl0OI
;
input
[
RABITS
:
0
]
CORETSE_AHBo0OI
;
input
[
RABITS
:
0
]
CORETSE_AHBi0OI
;
input
CORETSE_AHBO1OI
;
input
CORETSE_AHBI1OI
;
input
CORETSE_AHBIoo
;
input
[
RABITS
:
0
]
CORETSE_AHBiii
;
input
CORETSE_AHBIOOI
;
input
[
RABITS
:
0
]
CORETSE_AHBOOOI
;
output
CORETSE_AHBlIOI
;
output
CORETSE_AHBlIi
;
output
CORETSE_AHBoIi
;
output
CORETSE_AHBiIi
;
output
CORETSE_AHBlOOI
;
wire
CORETSE_AHBlIi
;
wire
CORETSE_AHBoIi
;
reg
CORETSE_AHBiIi
;
reg
CORETSE_AHBlOOI
;
parameter
CORETSE_AHBIoII
=
1
;
parameter
CORETSE_AHBoloI
=
{
RABITS
{
1
'b
0
}
}
;
parameter
CORETSE_AHBol0I
=
{
(
RABITS
+
1
)
{
1
'b
0
}
}
;
reg
[
5
:
0
]
CORETSE_AHBiOOl
;
reg
[
15
:
0
]
CORETSE_AHBOIOl
;
reg
[
6
:
0
]
CORETSE_AHBIIOl
;
reg
CORETSE_AHBlIOl
;
reg
CORETSE_AHBoIOl
;
wire
[
RABITS
:
0
]
CORETSE_AHBiIOl
;
reg
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBoooI
;
reg
[
RABITS
:
0
]
CORETSE_AHBiooI
;
reg
CORETSE_AHBOlOl
;
reg
CORETSE_AHBIlOl
;
reg
CORETSE_AHBllOl
;
reg
CORETSE_AHBolOl
;
reg
[
RABITS
:
0
]
CORETSE_AHBilOl
;
reg
[
RABITS
:
0
]
CORETSE_AHBO0Ol
;
reg
CORETSE_AHBI0Ol
;
reg
CORETSE_AHBl0Ol
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
01
;
else
if
(
CORETSE_AHBllo
)
case
(
CORETSE_AHBiOOl
)
6
'h
01
:
if
(
CORETSE_AHBlIOl
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
02
;
6
'h
02
:
if
(
~
CORETSE_AHBIoo
|
CORETSE_AHBI1OI
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
04
;
6
'h
04
:
if
(
CORETSE_AHBIoo
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
08
;
6
'h
08
:
if
(
~
CORETSE_AHBoIOl
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
10
;
else
if
(
~
(
|
CORETSE_AHBOIOl
)
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
02
;
6
'h
10
:
if
(
~
CORETSE_AHBIoo
|
CORETSE_AHBI1OI
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
20
;
6
'h
20
:
if
(
CORETSE_AHBIoo
)
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
01
;
default
:
CORETSE_AHBiOOl
<=
#
CORETSE_AHBIoII
6
'h
01
;
endcase
end
assign
CORETSE_AHBlIi
=
~
CORETSE_AHBI1OI
&
(
CORETSE_AHBiOOl
[
1
]
|
CORETSE_AHBiOOl
[
4
]
)
;
assign
CORETSE_AHBoIi
=
(
|
CORETSE_AHBiOOl
[
2
:
0
]
)
;
assign
CORETSE_AHBlIOI
=
~
CORETSE_AHBiOOl
[
0
]
|
CORETSE_AHBl0Ol
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBiIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBiIi
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1OI
&
(
CORETSE_AHBiOOl
[
1
]
|
(
CORETSE_AHBiIi
&
~
CORETSE_AHBiOOl
[
4
]
)
)
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBOIOl
<=
#
CORETSE_AHBIoII
16
'h
FFFF
;
else
if
(
CORETSE_AHBllo
)
begin
if
(
CORETSE_AHBiOOl
[
3
]
&
(
CORETSE_AHBOIOl
==
16
'h
0
)
)
CORETSE_AHBOIOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0OI
;
else
if
(
(
|
CORETSE_AHBiOOl
[
3
:
1
]
)
&
(
(
CORETSE_AHBO1OI
&
(
CORETSE_AHBIIOl
==
7
'd
126
)
)
|
(
~
CORETSE_AHBO1OI
&
(
CORETSE_AHBIIOl
==
7
'd
127
)
)
)
)
CORETSE_AHBOIOl
<=
#
CORETSE_AHBIoII
(
CORETSE_AHBOIOl
-
16
'h
1
)
;
else
if
(
~
(
|
CORETSE_AHBiOOl
[
3
:
1
]
)
)
CORETSE_AHBOIOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0OI
;
end
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBIIOl
<=
#
CORETSE_AHBIoII
7
'h
0
;
else
if
(
CORETSE_AHBllo
&
(
|
CORETSE_AHBiOOl
[
3
:
1
]
)
&
CORETSE_AHBO1OI
)
CORETSE_AHBIIOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIOl
+
7
'h
2
;
else
if
(
CORETSE_AHBllo
&
(
|
CORETSE_AHBiOOl
[
3
:
1
]
)
&
~
CORETSE_AHBO1OI
)
CORETSE_AHBIIOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIOl
+
7
'h
1
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBIIOl
<=
#
CORETSE_AHBIoII
7
'h
0
;
end
assign
CORETSE_AHBiIOl
=
(
~
CORETSE_AHBl0Ol
)
?
CORETSE_AHBol0I
:
(
CORETSE_AHBOlOl
==
CORETSE_AHBIlOl
)
?
{
1
'b
0
,
CORETSE_AHBoooI
}
:
CORETSE_AHBiooI
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBlIOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBlIOl
<=
#
CORETSE_AHBIoII
(
CORETSE_AHBiIOl
>
CORETSE_AHBo0OI
)
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBoIOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBoIOl
<=
#
CORETSE_AHBIoII
(
CORETSE_AHBiIOl
>
CORETSE_AHBi0OI
)
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBoooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoloI
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBoooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBilOl
[
(
RABITS
-
1
)
:
0
]
-
CORETSE_AHBO0Ol
[
(
RABITS
-
1
)
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBiooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBiooI
<=
#
CORETSE_AHBIoII
{
1
'b
1
,
CORETSE_AHBilOl
[
(
RABITS
-
1
)
:
0
]
}
-
{
1
'b
0
,
CORETSE_AHBO0Ol
[
(
RABITS
-
1
)
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBOlOl
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBOlOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBilOl
[
RABITS
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBIlOl
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBIlOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0Ol
[
RABITS
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBllOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBllOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOOI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBolOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBolOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBllOl
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBlOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBlOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBolOl
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBilOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBolOl
&
~
CORETSE_AHBlOOI
)
CORETSE_AHBilOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBiii
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBO0Ol
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBolOl
&
~
CORETSE_AHBlOOI
)
CORETSE_AHBO0Ol
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOOI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBI0Ol
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI0Ol
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOII
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBo0II
)
begin
if
(
CORETSE_AHBo0II
)
CORETSE_AHBl0Ol
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl0Ol
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0Ol
;
end
endmodule
