// REVISION    : $Revision: 1.4 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
perex_pcs
#
(
parameter
CORETSE_AHBlOI
=
1
'b
0
)
(
CORETSE_AHBOO1
,
CORETSE_AHBiO11
,
CORETSE_AHBOI11
,
CORETSE_AHBl01
,
CORETSE_AHBoii0
,
CORETSE_AHBioO1
,
CORETSE_AHBlO11
,
CORETSE_AHBOO11
,
CORETSE_AHBlo01
,
CORETSE_AHBi010
,
CORETSE_AHBiIO1
,
CORETSE_AHBOo1
,
CORETSE_AHBOIO1
,
CORETSE_AHBIIO1
,
CORETSE_AHBlIO1
,
CORETSE_AHBoIO1
,
CORETSE_AHBIii0
,
CORETSE_AHBOii0
,
CORETSE_AHBlii0
)
;
input
CORETSE_AHBOO1
;
input
[
19
:
0
]
CORETSE_AHBiO11
;
input
CORETSE_AHBOI11
;
input
CORETSE_AHBl01
;
input
CORETSE_AHBoii0
;
input
[
1
:
0
]
CORETSE_AHBioO1
;
input
CORETSE_AHBlO11
;
input
CORETSE_AHBOO11
;
input
CORETSE_AHBlo01
;
input
CORETSE_AHBi010
;
input
CORETSE_AHBiIO1
;
output
CORETSE_AHBOo1
;
output
CORETSE_AHBOIO1
;
output
CORETSE_AHBIIO1
;
output
CORETSE_AHBlIO1
;
output
[
15
:
0
]
CORETSE_AHBoIO1
;
output
[
1
:
0
]
CORETSE_AHBIii0
;
output
[
15
:
0
]
CORETSE_AHBOii0
;
output
[
1
:
0
]
CORETSE_AHBlii0
;
reg
CORETSE_AHBOo1
;
wire
CORETSE_AHBOIO1
;
wire
CORETSE_AHBIIO1
;
reg
CORETSE_AHBlIO1
;
reg
[
15
:
0
]
CORETSE_AHBoIO1
;
reg
[
1
:
0
]
CORETSE_AHBIii0
;
reg
[
15
:
0
]
CORETSE_AHBOii0
;
reg
[
1
:
0
]
CORETSE_AHBlii0
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBiOoi
,
CORETSE_AHBOIoi
,
CORETSE_AHBIIoi
,
CORETSE_AHBlIoi
;
reg
[
1
:
0
]
CORETSE_AHBoIoi
,
CORETSE_AHBiIoi
;
wire
[
1
:
0
]
CORETSE_AHBOloi
;
wire
CORETSE_AHBIloi
;
reg
CORETSE_AHBlloi
;
wire
[
15
:
0
]
CORETSE_AHBoloi
;
wire
[
5
:
0
]
CORETSE_AHBiloi
;
wire
[
1
:
0
]
CORETSE_AHBO0oi
;
wire
[
1
:
0
]
CORETSE_AHBI0oi
;
reg
[
31
:
0
]
CORETSE_AHBl0oi
;
reg
[
11
:
0
]
CORETSE_AHBo0oi
;
reg
[
3
:
0
]
CORETSE_AHBi0oi
;
wire
CORETSE_AHBO1oi
;
wire
[
7
:
0
]
CORETSE_AHBI1oi
;
wire
CORETSE_AHBl1oi
,
CORETSE_AHBo1oi
,
CORETSE_AHBi1oi
,
CORETSE_AHBOooi
;
wire
CORETSE_AHBIooi
,
CORETSE_AHBlooi
;
wire
CORETSE_AHBoooi
;
wire
CORETSE_AHBiooi
;
wire
CORETSE_AHBOioi
,
CORETSE_AHBIioi
;
wire
CORETSE_AHBlioi
,
CORETSE_AHBoioi
;
wire
CORETSE_AHBiioi
,
CORETSE_AHBOOii
;
wire
CORETSE_AHBIOii
;
wire
CORETSE_AHBlOii
,
CORETSE_AHBoOii
;
wire
CORETSE_AHBiOii
;
wire
CORETSE_AHBOIii
,
CORETSE_AHBIIii
;
wire
CORETSE_AHBlIii
,
CORETSE_AHBoIii
;
wire
CORETSE_AHBiIii
,
CORETSE_AHBOlii
;
wire
CORETSE_AHBIlii
,
CORETSE_AHBllii
;
wire
CORETSE_AHBolii
;
wire
CORETSE_AHBilii
;
wire
CORETSE_AHBO0ii
,
CORETSE_AHBI0ii
;
wire
CORETSE_AHBl0ii
;
wire
CORETSE_AHBo0ii
;
wire
CORETSE_AHBi0ii
;
wire
CORETSE_AHBO1ii
;
wire
CORETSE_AHBI1ii
;
wire
CORETSE_AHBl1ii
,
CORETSE_AHBo1ii
;
wire
[
1
:
0
]
CORETSE_AHBi1ii
;
reg
[
1
:
0
]
CORETSE_AHBOoii
;
wire
CORETSE_AHBIoii
,
CORETSE_AHBloii
,
CORETSE_AHBooii
;
wire
CORETSE_AHBioii
;
wire
CORETSE_AHBOiii
;
reg
CORETSE_AHBIiii
;
wire
CORETSE_AHBliii
,
CORETSE_AHBoiii
;
reg
CORETSE_AHBiiii
,
CORETSE_AHBOOOOI
;
wire
CORETSE_AHBIOOOI
;
reg
CORETSE_AHBlOOOI
;
wire
CORETSE_AHBoOOOI
,
CORETSE_AHBiOOOI
;
wire
CORETSE_AHBOIOOI
,
CORETSE_AHBIIOOI
;
wire
CORETSE_AHBlIOOI
,
CORETSE_AHBoIOOI
;
reg
CORETSE_AHBiIOOI
,
CORETSE_AHBOlOOI
;
reg
CORETSE_AHBIlOOI
,
CORETSE_AHBllOOI
;
reg
CORETSE_AHBolOOI
,
CORETSE_AHBilOOI
;
wire
CORETSE_AHBO0OOI
;
wire
CORETSE_AHBI0OOI
,
CORETSE_AHBl0OOI
,
CORETSE_AHBo0OOI
,
CORETSE_AHBi0OOI
;
wire
CORETSE_AHBO1OOI
;
reg
CORETSE_AHBI1OOI
;
wire
CORETSE_AHBl1OOI
;
reg
CORETSE_AHBo1OOI
;
wire
CORETSE_AHBi1OOI
;
reg
CORETSE_AHBOoOOI
;
wire
CORETSE_AHBIoOOI
;
reg
CORETSE_AHBloOOI
;
wire
CORETSE_AHBooOOI
;
reg
CORETSE_AHBioOOI
;
wire
CORETSE_AHBOiOOI
;
reg
CORETSE_AHBIiOOI
;
wire
CORETSE_AHBliOOI
;
reg
CORETSE_AHBoiOOI
;
wire
CORETSE_AHBiiOOI
;
wire
[
15
:
0
]
CORETSE_AHBOOIOI
;
wire
CORETSE_AHBIOIOI
;
reg
CORETSE_AHBlOIOI
;
reg
CORETSE_AHBoOIOI
;
wire
CORETSE_AHBiOIOI
;
reg
CORETSE_AHBOIIOI
;
wire
CORETSE_AHBIIIOI
;
reg
CORETSE_AHBlIIOI
;
wire
CORETSE_AHBoIIOI
;
reg
CORETSE_AHBiIIOI
;
wire
CORETSE_AHBOlIOI
;
reg
CORETSE_AHBIlIOI
;
wire
CORETSE_AHBllIOI
;
reg
CORETSE_AHBolIOI
;
wire
CORETSE_AHBilIOI
;
reg
CORETSE_AHBO0IOI
;
wire
CORETSE_AHBI0IOI
;
reg
CORETSE_AHBl0IOI
;
wire
[
1
:
0
]
CORETSE_AHBo0IOI
;
wire
[
1
:
0
]
CORETSE_AHBi0IOI
,
CORETSE_AHBO1IOI
;
wire
[
15
:
0
]
CORETSE_AHBI1IOI
;
reg
CORETSE_AHBl1IOI
;
reg
CORETSE_AHBo1IOI
;
assign
CORETSE_AHBi1IOI
=
1
'b
0
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiOoi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiOoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBl01
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOIoi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOIoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOoi
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIIoi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIIoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIoi
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlIoi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlIoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIoi
^
CORETSE_AHBIIoi
|
CORETSE_AHBOI11
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoIoi
[
1
:
0
]
<=
#
CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBoIoi
[
1
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBioO1
[
1
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiIoi
[
1
:
0
]
<=
#
CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBiIoi
[
1
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIoi
[
1
:
0
]
;
end
assign
CORETSE_AHBOloi
[
0
]
=
~
CORETSE_AHBOO11
&
CORETSE_AHBlloi
;
assign
CORETSE_AHBOloi
[
1
]
=
~
CORETSE_AHBOO11
&
CORETSE_AHBO0oi
[
0
]
;
assign
CORETSE_AHBIloi
=
~
CORETSE_AHBOO11
&
CORETSE_AHBO0oi
[
1
]
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlloi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlloi
<=
#
CORETSE_AHBIoII
CORETSE_AHBIloi
;
end
r10b8b
CORETSE_AHBOoIOI
(
.CORETSE_AHBIoIOI
(
CORETSE_AHBiO11
[
9
:
0
]
)
,
.CORETSE_AHBOloi
(
CORETSE_AHBOloi
[
0
]
)
,
.CORETSE_AHBOo1
(
CORETSE_AHBOo1
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBI1oi
[
7
:
0
]
)
,
.CORETSE_AHBo0oi
(
CORETSE_AHBiloi
[
2
:
0
]
)
,
.CORETSE_AHBO0oi
(
CORETSE_AHBO0oi
[
0
]
)
,
.CORETSE_AHBi0oi
(
CORETSE_AHBI0oi
[
0
]
)
)
;
r10b8b
CORETSE_AHBloIOI
(
.CORETSE_AHBIoIOI
(
CORETSE_AHBiO11
[
19
:
10
]
)
,
.CORETSE_AHBOloi
(
CORETSE_AHBOloi
[
1
]
)
,
.CORETSE_AHBOo1
(
CORETSE_AHBOo1
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBoloi
[
15
:
8
]
)
,
.CORETSE_AHBo0oi
(
CORETSE_AHBiloi
[
5
:
3
]
)
,
.CORETSE_AHBO0oi
(
CORETSE_AHBO0oi
[
1
]
)
,
.CORETSE_AHBi0oi
(
CORETSE_AHBI0oi
[
1
]
)
)
;
assign
CORETSE_AHBO1oi
=
(
CORETSE_AHBiO11
[
9
:
0
]
==
10
'h
27c
)
|
(
CORETSE_AHBiO11
[
9
:
0
]
==
10
'h
183
)
;
assign
CORETSE_AHBoloi
[
7
:
0
]
=
(
{
8
{
CORETSE_AHBO1oi
}
}
&
8
'h
3c
)
|
(
{
8
{
~
CORETSE_AHBO1oi
}
}
&
CORETSE_AHBI1oi
[
7
:
0
]
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBl0oi
[
31
:
0
]
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
CORETSE_AHBl0oi
[
31
:
0
]
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBoloi
[
15
:
0
]
,
CORETSE_AHBl0oi
[
31
:
16
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBo0oi
[
11
:
0
]
<=
#
CORETSE_AHBIoII
12
'h
0
;
else
CORETSE_AHBo0oi
[
11
:
0
]
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBiloi
[
5
:
0
]
,
CORETSE_AHBo0oi
[
11
:
6
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBi0oi
[
3
:
0
]
<=
#
CORETSE_AHBIoII
4
'h
0
;
else
CORETSE_AHBi0oi
[
3
:
0
]
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBI0oi
[
1
:
0
]
,
CORETSE_AHBi0oi
[
3
:
2
]
}
;
end
assign
CORETSE_AHBl1oi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
000
;
assign
CORETSE_AHBo1oi
=
CORETSE_AHBo0oi
[
2
:
0
]
!=
3
'b
000
;
assign
CORETSE_AHBIooi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
001
;
assign
CORETSE_AHBlooi
=
CORETSE_AHBo0oi
[
2
:
0
]
!=
3
'b
001
;
assign
CORETSE_AHBoooi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
010
;
assign
CORETSE_AHBiooi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
011
;
assign
CORETSE_AHBOioi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
100
;
assign
CORETSE_AHBIioi
=
CORETSE_AHBo0oi
[
2
:
0
]
!=
3
'b
100
;
assign
CORETSE_AHBlioi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
100
&
CORETSE_AHBl0oi
[
7
:
0
]
==
8
'h
BC
;
assign
CORETSE_AHBoioi
=
CORETSE_AHBo0oi
[
2
:
0
]
!=
3
'b
100
|
CORETSE_AHBl0oi
[
7
:
0
]
!=
8
'h
BC
;
assign
CORETSE_AHBiioi
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
101
;
assign
CORETSE_AHBOOii
=
CORETSE_AHBo0oi
[
2
:
0
]
!=
3
'b
101
;
assign
CORETSE_AHBIOii
=
CORETSE_AHBo0oi
[
2
:
0
]
==
3
'b
111
;
assign
CORETSE_AHBlOii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
001
;
assign
CORETSE_AHBoOii
=
CORETSE_AHBo0oi
[
5
:
3
]
!=
3
'b
001
;
assign
CORETSE_AHBiOii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
010
;
assign
CORETSE_AHBOIii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
011
;
assign
CORETSE_AHBIIii
=
CORETSE_AHBo0oi
[
5
:
3
]
!=
3
'b
011
;
assign
CORETSE_AHBlIii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
100
;
assign
CORETSE_AHBoIii
=
CORETSE_AHBo0oi
[
5
:
3
]
!=
3
'b
100
;
assign
CORETSE_AHBiIii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
100
&
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
BC
;
assign
CORETSE_AHBOlii
=
CORETSE_AHBo0oi
[
5
:
3
]
!=
3
'b
100
|
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
BC
;
assign
CORETSE_AHBIlii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
101
;
assign
CORETSE_AHBllii
=
CORETSE_AHBo0oi
[
5
:
3
]
!=
3
'b
101
;
assign
CORETSE_AHBolii
=
CORETSE_AHBo0oi
[
5
:
3
]
==
3
'b
111
;
assign
CORETSE_AHBi1oi
=
CORETSE_AHBo0oi
[
8
:
6
]
==
3
'b
000
;
assign
CORETSE_AHBilii
=
CORETSE_AHBo0oi
[
8
:
6
]
==
3
'b
001
;
assign
CORETSE_AHBO0ii
=
CORETSE_AHBo0oi
[
8
:
6
]
==
3
'b
011
;
assign
CORETSE_AHBI0ii
=
CORETSE_AHBo0oi
[
8
:
6
]
!=
3
'b
011
;
assign
CORETSE_AHBl0ii
=
CORETSE_AHBo0oi
[
8
:
6
]
==
3
'b
100
&
CORETSE_AHBl0oi
[
23
:
16
]
==
8
'h
BC
;
assign
CORETSE_AHBo0ii
=
CORETSE_AHBo0oi
[
8
:
6
]
==
3
'b
101
;
assign
CORETSE_AHBi0ii
=
CORETSE_AHBo0oi
[
11
:
9
]
==
3
'b
001
;
assign
CORETSE_AHBO1ii
=
CORETSE_AHBo0oi
[
11
:
9
]
==
3
'b
011
;
assign
CORETSE_AHBI1ii
=
CORETSE_AHBo0oi
[
11
:
9
]
==
3
'b
100
&
CORETSE_AHBl0oi
[
31
:
24
]
==
8
'h
BC
;
assign
CORETSE_AHBOooi
=
CORETSE_AHBo0oi
[
11
:
9
]
==
3
'b
000
;
assign
CORETSE_AHBl1ii
=
CORETSE_AHBIooi
;
assign
CORETSE_AHBo1ii
=
~
CORETSE_AHBl1ii
;
assign
CORETSE_AHBi1ii
=
{
2
{
CORETSE_AHBlOOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBiIOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
10
|
{
2
{
CORETSE_AHBiIOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBIlOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
10
|
{
2
{
CORETSE_AHBIlOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBolOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
10
|
{
2
{
CORETSE_AHBOlOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBIoii
}
}
&
2
'b
11
|
{
2
{
CORETSE_AHBOlOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBIoii
}
}
&
2
'b
11
|
{
2
{
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBooii
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBllOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBilOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBIoii
}
}
&
2
'b
11
|
{
2
{
CORETSE_AHBilOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBooii
}
}
&
2
'b
01
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOoii
<=
#
CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBOoii
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1ii
;
end
assign
CORETSE_AHBIoii
=
CORETSE_AHBOoii
==
2
'b
01
;
assign
CORETSE_AHBloii
=
CORETSE_AHBOoii
==
2
'b
10
;
assign
CORETSE_AHBooii
=
CORETSE_AHBOoii
==
2
'b
11
;
assign
CORETSE_AHBioii
=
CORETSE_AHBoii0
|
CORETSE_AHBlo01
;
assign
CORETSE_AHBOiii
=
CORETSE_AHBlIoi
&
~
CORETSE_AHBioii
|
CORETSE_AHBIiii
&
(
~
CORETSE_AHBOIoi
&
~
CORETSE_AHBioii
|
CORETSE_AHBIioi
|
CORETSE_AHBllii
)
|
CORETSE_AHBiiii
&
(
CORETSE_AHBIooi
|
CORETSE_AHBlOii
|
CORETSE_AHBlIii
|
CORETSE_AHBOioi
&
CORETSE_AHBllii
)
|
CORETSE_AHBOOOOI
&
(
CORETSE_AHBIooi
|
CORETSE_AHBlOii
|
CORETSE_AHBlIii
|
CORETSE_AHBOioi
&
CORETSE_AHBllii
)
|
CORETSE_AHBIlOOI
&
CORETSE_AHBIooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBllOOI
&
CORETSE_AHBIooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBolOOI
&
(
CORETSE_AHBIooi
|
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBilOOI
&
(
CORETSE_AHBIooi
|
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
&
(
CORETSE_AHBIoii
|
CORETSE_AHBloii
)
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIiii
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBIiii
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiii
;
end
assign
CORETSE_AHBliii
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBIiii
&
CORETSE_AHBOioi
&
CORETSE_AHBIlii
|
CORETSE_AHBiiii
&
CORETSE_AHBIioi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiiii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiiii
<=
#
CORETSE_AHBIoII
CORETSE_AHBliii
;
end
assign
CORETSE_AHBoiii
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBiiii
&
CORETSE_AHBOioi
&
CORETSE_AHBIlii
|
CORETSE_AHBOOOOI
&
CORETSE_AHBIioi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOOOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOOOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiii
;
end
assign
CORETSE_AHBIOOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBOOOOI
&
CORETSE_AHBOioi
&
CORETSE_AHBIlii
|
CORETSE_AHBlOOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBOlOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
(
CORETSE_AHBloii
|
CORETSE_AHBooii
)
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlOOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlOOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOOOI
;
end
assign
CORETSE_AHBoOOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBlOOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBOlOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
&
CORETSE_AHBooii
|
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBloii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiIOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiIOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOOOI
;
end
assign
CORETSE_AHBiOOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBlOOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBiIOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBOlOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBIoii
|
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBooii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOlOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOlOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOOOI
;
end
assign
CORETSE_AHBOIOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBlOOOI
&
CORETSE_AHBIooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBiIOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBOlOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
&
(
CORETSE_AHBIoii
|
CORETSE_AHBloii
)
|
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
&
CORETSE_AHBooii
|
CORETSE_AHBilOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBloii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIlOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIlOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIOOI
;
end
assign
CORETSE_AHBIIOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBiIOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBOlOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBIlOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBIoii
|
CORETSE_AHBilOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBooii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBllOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBllOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIOOI
;
end
assign
CORETSE_AHBlIOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBiIOOI
&
CORETSE_AHBIooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBOlOOI
&
CORETSE_AHBIooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBIlOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
|
CORETSE_AHBllOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
&
(
CORETSE_AHBIoii
|
CORETSE_AHBloii
)
|
CORETSE_AHBilOOI
&
CORETSE_AHBlooi
&
(
CORETSE_AHBlOii
|
CORETSE_AHBlIii
)
&
CORETSE_AHBooii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBolOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBolOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIOOI
;
end
assign
CORETSE_AHBoIOOI
=
(
CORETSE_AHBOIoi
&
~
CORETSE_AHBlIoi
|
CORETSE_AHBioii
)
&
(
CORETSE_AHBIlOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBllOOI
&
CORETSE_AHBIooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBolOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
|
CORETSE_AHBilOOI
&
CORETSE_AHBlooi
&
CORETSE_AHBoOii
&
CORETSE_AHBoIii
&
CORETSE_AHBIoii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBilOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBilOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIOOI
;
end
assign
CORETSE_AHBO0OOI
=
~
CORETSE_AHBOo1
&
CORETSE_AHBIOOOI
|
CORETSE_AHBOo1
&
~
CORETSE_AHBOiii
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOo1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0OOI
;
end
assign
CORETSE_AHBI0OOI
=
CORETSE_AHBiIoi
[
1
:
0
]
==
2
'b
00
;
assign
CORETSE_AHBl0OOI
=
CORETSE_AHBiIoi
[
1
:
0
]
==
2
'b
01
;
assign
CORETSE_AHBo0OOI
=
(
CORETSE_AHBiIoi
[
1
:
0
]
==
2
'b
10
)
|
~
CORETSE_AHBo1IOI
;
assign
CORETSE_AHBi0OOI
=
~
CORETSE_AHBo0OOI
;
assign
CORETSE_AHBO1OOI
=
~
CORETSE_AHBI1OOI
&
~
CORETSE_AHBO0OOI
|
CORETSE_AHBI1OOI
&
~
CORETSE_AHBO0OOI
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBI1OOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI1OOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1OOI
;
end
assign
CORETSE_AHBl1OOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBI1OOI
&
CORETSE_AHBoioi
|
CORETSE_AHBoiOOI
&
CORETSE_AHBoioi
|
CORETSE_AHBo1OOI
&
CORETSE_AHBoioi
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBo1OOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBo1OOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1OOI
;
end
assign
CORETSE_AHBi1OOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBi0OOI
&
CORETSE_AHBlioi
&
CORETSE_AHBIlii
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
B5
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
42
|
CORETSE_AHBo0OOI
&
CORETSE_AHBlioi
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
B5
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
42
|
CORETSE_AHBOoOOI
&
CORETSE_AHBi0OOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBIlii
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
B5
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
42
|
CORETSE_AHBOoOOI
&
CORETSE_AHBo0OOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
B5
&
CORETSE_AHBl0oi
[
15
:
8
]
!=
8
'h
42
|
CORETSE_AHBloOOI
&
CORETSE_AHBlioi
|
CORETSE_AHBIlIOI
&
CORETSE_AHBlioi
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOoOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOoOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1OOI
;
end
assign
CORETSE_AHBOIO1
=
CORETSE_AHBOoOOI
;
assign
CORETSE_AHBooOOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBo1OOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBIlii
&
(
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
B5
|
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
42
)
|
CORETSE_AHBOoOOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBIlii
&
(
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
B5
|
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
42
)
|
CORETSE_AHBIiOOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBIlii
&
(
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
B5
|
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
42
)
|
CORETSE_AHBoiOOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBIlii
&
(
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
B5
|
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
42
)
|
CORETSE_AHBolIOI
&
(
CORETSE_AHBlioi
|
CORETSE_AHBi0oi
[
0
]
)
&
CORETSE_AHBIlii
&
(
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
B5
|
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
42
)
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBioOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBioOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBooOOI
;
end
assign
CORETSE_AHBOiOOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBioOOI
&
CORETSE_AHBiioi
&
CORETSE_AHBIlii
|
CORETSE_AHBIlIOI
&
CORETSE_AHBiioi
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIiOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIiOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiOOI
;
end
assign
CORETSE_AHBiiOOI
=
CORETSE_AHBOiOOI
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlIO1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlIO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiOOI
;
end
assign
CORETSE_AHBOOIOI
[
15
:
0
]
=
{
16
{
CORETSE_AHBOiOOI
}
}
&
{
CORETSE_AHBl0oi
[
15
:
0
]
}
|
{
16
{
~
CORETSE_AHBOiOOI
}
}
&
{
CORETSE_AHBoIO1
[
15
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoIO1
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBoIO1
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOIOI
[
15
:
0
]
;
end
assign
CORETSE_AHBliOOI
=
CORETSE_AHBI1OOI
|
CORETSE_AHBOo1
&
(
CORETSE_AHBOoOOI
&
CORETSE_AHBi0OOI
&
(
CORETSE_AHBoioi
|
CORETSE_AHBllii
|
CORETSE_AHBOI11
)
|
CORETSE_AHBioOOI
&
(
CORETSE_AHBOOii
|
CORETSE_AHBllii
|
CORETSE_AHBOI11
)
|
CORETSE_AHBIiOOI
&
(
CORETSE_AHBoioi
|
CORETSE_AHBIooi
|
CORETSE_AHBlOii
)
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoiOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoiOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBliOOI
;
end
assign
CORETSE_AHBIIO1
=
CORETSE_AHBoiOOI
;
assign
CORETSE_AHBIoOOI
=
CORETSE_AHBOoOOI
&
CORETSE_AHBo0OOI
&
CORETSE_AHBoioi
&
~
CORETSE_AHBi0oi
[
0
]
&
CORETSE_AHBo1oi
|
CORETSE_AHBloOOI
&
CORETSE_AHBoioi
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBloOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBloOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoOOI
;
end
assign
CORETSE_AHBIOIOI
=
(
CORETSE_AHBOoOOI
&
CORETSE_AHBo0OOI
&
CORETSE_AHBoioi
&
~
CORETSE_AHBi0oi
[
0
]
&
CORETSE_AHBl1oi
)
|
CORETSE_AHBoOIOI
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlOIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlOIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOIOI
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoOIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoOIOI
<=
#
CORETSE_AHBIoII
(
CORETSE_AHBO0IOI
&
(
(
CORETSE_AHBiooi
&
CORETSE_AHBOIii
&
CORETSE_AHBi1oi
)
|
(
CORETSE_AHBOIii
&
CORETSE_AHBO0ii
&
CORETSE_AHBOooi
)
)
)
;
end
assign
CORETSE_AHBiOIOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBIOIOI
|
CORETSE_AHBOIIOI
&
(
CORETSE_AHBIIIOI
|
CORETSE_AHBoIIOI
)
&
~
CORETSE_AHBI0IOI
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOIIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOIIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOIOI
;
end
assign
CORETSE_AHBIIIOI
=
CORETSE_AHBOo1
&
CORETSE_AHBOIIOI
&
CORETSE_AHBiioi
&
CORETSE_AHBIlii
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlIIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlIIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIIOI
;
end
assign
CORETSE_AHBoIIOI
=
CORETSE_AHBOo1
&
CORETSE_AHBOIIOI
&
(
~
CORETSE_AHBIIIOI
&
~
CORETSE_AHBOlIOI
&
~
CORETSE_AHBllIOI
&
~
CORETSE_AHBilIOI
|
CORETSE_AHBIOii
|
CORETSE_AHBolii
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiIIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiIIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIIOI
;
end
assign
CORETSE_AHBOlIOI
=
CORETSE_AHBOo1
&
CORETSE_AHBOIIOI
&
(
CORETSE_AHBlioi
&
CORETSE_AHBIlii
&
CORETSE_AHBl0ii
|
CORETSE_AHBlioi
&
CORETSE_AHBIlii
&
(
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
B5
|
CORETSE_AHBl0oi
[
15
:
8
]
==
8
'h
42
)
&
CORETSE_AHBo0ii
&
CORETSE_AHBl0oi
[
23
:
16
]
==
8
'h
00
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIlIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIlIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOlIOI
;
end
assign
CORETSE_AHBllIOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBOIIOI
&
CORETSE_AHBoooi
&
CORETSE_AHBOIii
&
CORETSE_AHBl0ii
|
CORETSE_AHBO0IOI
&
CORETSE_AHBiooi
&
CORETSE_AHBOIii
&
CORETSE_AHBl0ii
|
CORETSE_AHBolIOI
&
CORETSE_AHBoioi
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBolIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBolIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBllIOI
;
end
assign
CORETSE_AHBilIOI
=
CORETSE_AHBOo1
&
(
(
CORETSE_AHBOIIOI
&
CORETSE_AHBiOii
&
CORETSE_AHBO0ii
&
CORETSE_AHBO1ii
)
|
(
CORETSE_AHBOIIOI
&
CORETSE_AHBoooi
&
CORETSE_AHBOIii
&
CORETSE_AHBO0ii
)
|
(
CORETSE_AHBO0IOI
&
CORETSE_AHBiooi
&
CORETSE_AHBOIii
&
CORETSE_AHBO0ii
)
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBO0IOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO0IOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBilIOI
;
end
assign
CORETSE_AHBI0IOI
=
CORETSE_AHBOo1
&
(
CORETSE_AHBOIIOI
&
CORETSE_AHBiooi
&
CORETSE_AHBOIii
&
CORETSE_AHBO0ii
)
|
(
CORETSE_AHBOIIOI
&
CORETSE_AHBOIii
&
CORETSE_AHBO0ii
&
CORETSE_AHBO1ii
&
~
CORETSE_AHBoooi
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBl0IOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl0IOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0IOI
;
end
assign
CORETSE_AHBi0IOI
[
1
]
=
CORETSE_AHBIoOOI
|
CORETSE_AHBoIIOI
&
CORETSE_AHBolii
|
CORETSE_AHBoIIOI
&
CORETSE_AHBi0ii
|
CORETSE_AHBoIIOI
&
CORETSE_AHBiOii
&
CORETSE_AHBO0ii
&
CORETSE_AHBI1ii
|
CORETSE_AHBoIIOI
&
CORETSE_AHBiOii
&
CORETSE_AHBI0ii
&
CORETSE_AHBO1ii
|
CORETSE_AHBoIIOI
&
CORETSE_AHBoooi
&
CORETSE_AHBIIii
&
CORETSE_AHBl0ii
|
CORETSE_AHBilIOI
;
assign
CORETSE_AHBi0IOI
[
0
]
=
CORETSE_AHBIoOOI
|
CORETSE_AHBoIIOI
&
CORETSE_AHBIOii
|
CORETSE_AHBoIIOI
&
CORETSE_AHBilii
|
CORETSE_AHBoIIOI
&
CORETSE_AHBiOii
&
CORETSE_AHBO0ii
&
CORETSE_AHBI1ii
|
CORETSE_AHBOlIOI
&
~
CORETSE_AHBIlIOI
|
CORETSE_AHBilIOI
&
CORETSE_AHBoooi
|
CORETSE_AHBO0IOI
&
CORETSE_AHBilIOI
|
CORETSE_AHBI0IOI
;
assign
CORETSE_AHBO1IOI
[
1
]
=
~
CORETSE_AHBlO11
&
CORETSE_AHBi0IOI
[
1
]
|
CORETSE_AHBlO11
&
CORETSE_AHBiO11
[
19
]
;
assign
CORETSE_AHBO1IOI
[
0
]
=
~
CORETSE_AHBlO11
&
CORETSE_AHBi0IOI
[
0
]
|
CORETSE_AHBlO11
&
CORETSE_AHBiO11
[
9
]
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlii0
[
1
:
0
]
<=
#
CORETSE_AHBIoII
2
'b
0
;
else
CORETSE_AHBlii0
[
1
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1IOI
[
1
:
0
]
;
end
assign
CORETSE_AHBo0IOI
[
1
]
=
~
CORETSE_AHBlO11
&
(
CORETSE_AHBIOIOI
|
CORETSE_AHBIii0
[
0
]
&
~
(
CORETSE_AHBl1OOI
|
CORETSE_AHBi1OOI
|
CORETSE_AHBooOOI
|
CORETSE_AHBOiOOI
|
CORETSE_AHBllIOI
|
CORETSE_AHBilIOI
|
CORETSE_AHBl0IOI
)
)
|
CORETSE_AHBlO11
&
CORETSE_AHBiO11
[
18
]
;
assign
CORETSE_AHBo0IOI
[
0
]
=
~
CORETSE_AHBlO11
&
(
CORETSE_AHBIOIOI
|
CORETSE_AHBIii0
[
0
]
&
~
(
CORETSE_AHBl1OOI
|
CORETSE_AHBi1OOI
&
~
(
CORETSE_AHBOlIOI
&
~
CORETSE_AHBIlIOI
)
|
CORETSE_AHBooOOI
|
CORETSE_AHBOiOOI
|
(
CORETSE_AHBilIOI
&
CORETSE_AHBoooi
)
|
(
CORETSE_AHBilIOI
&
CORETSE_AHBO0IOI
)
|
CORETSE_AHBllIOI
|
CORETSE_AHBl0IOI
)
)
|
CORETSE_AHBlO11
&
CORETSE_AHBiO11
[
8
]
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIii0
[
1
:
0
]
<=
#
CORETSE_AHBIoII
2
'b
0
;
else
CORETSE_AHBIii0
[
1
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0IOI
[
1
:
0
]
;
end
assign
CORETSE_AHBI1IOI
[
15
:
0
]
=
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBIoOOI
}
}
&
16
'h
0E0E
|
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBIOIOI
}
}
&
16
'h
5555
|
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBIIIOI
}
}
&
CORETSE_AHBl0oi
[
15
:
0
]
|
{
{
8
{
~
CORETSE_AHBlO11
&
CORETSE_AHBOIIOI
&
CORETSE_AHBoIIOI
&
~
CORETSE_AHBi0IOI
[
1
]
}
}
&
CORETSE_AHBl0oi
[
15
:
8
]
,
{
8
{
~
CORETSE_AHBlO11
&
CORETSE_AHBOIIOI
&
CORETSE_AHBoIIOI
&
~
CORETSE_AHBi0IOI
[
0
]
}
}
&
CORETSE_AHBl0oi
[
7
:
0
]
}
|
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBilIOI
&
CORETSE_AHBiOii
}
}
&
{
8
'h
0F
,
CORETSE_AHBl0oi
[
7
:
0
]
}
|
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBilIOI
&
CORETSE_AHBoooi
}
}
&
{
8
'h
0F
,
8
'h
0F
}
|
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBilIOI
&
~
CORETSE_AHBiOii
&
~
CORETSE_AHBoooi
}
}
&
{
8
'h
0F
,
8
'h
0F
}
|
{
16
{
~
CORETSE_AHBlO11
&
CORETSE_AHBO0IOI
&
CORETSE_AHBiooi
&
CORETSE_AHBOIii
&
CORETSE_AHBi1oi
}
}
&
{
8
'h
0F
,
8
'h
0F
}
|
{
16
{
CORETSE_AHBlO11
}
}
&
{
CORETSE_AHBiO11
[
17
:
10
]
,
CORETSE_AHBiO11
[
7
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOii0
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBOii0
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1IOI
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBl1IOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1IOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIO1
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBo1IOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo1IOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1IOI
;
end
endmodule
