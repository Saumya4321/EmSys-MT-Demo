//                     Proprietary and Confidential
// REVISION : $Revision: $
`include "include.v"
module
ptp_rtc
#
(
parameter
CORETSE_AHBlII
=
2
,
parameter
CORETSE_AHBIII
=
1
,
parameter
CORETSE_AHBiII
=
2
,
parameter
CORETSE_AHBoII
=
1
)
(
input
CORETSE_AHBIl0,
input
CORETSE_AHBOl0,
input
CORETSE_AHBOo0lI,
input
CORETSE_AHBl0I,
input
CORETSE_AHBlOo0I,
input
[
7
:
0
]
CORETSE_AHBolO1I,
input
[
7
:
0
]
CORETSE_AHBilO1I,
input
CORETSE_AHBO0O1I,
input
CORETSE_AHBI0O1I,
input
[
79
:
0
]
CORETSE_AHBl0O1I,
input
[
79
:
0
]
CORETSE_AHBo0O1I,
input
CORETSE_AHBoOo0I,
input
CORETSE_AHBi0O1I,
input
CORETSE_AHBO1O1I,
input
[
79
:
0
]
CORETSE_AHBI1O1I,
input
CORETSE_AHBl1O1I,
input
CORETSE_AHBo1O1I,
input
CORETSE_AHBi1O1I,
input
CORETSE_AHBOoO1I,
input
CORETSE_AHBIoO1I,
input
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
CORETSE_AHBloO1I,
input
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
CORETSE_AHBooO1I,
input
CORETSE_AHBioO1I,
input
[
`CORETSE_AHBIoI0
:
0
]
CORETSE_AHBOiO1I,
input
CORETSE_AHBIiO1I,
output
CORETSE_AHBliO1I,
output
CORETSE_AHBll0,
output
CORETSE_AHBoiO1I,
output
[
79
:
0
]
CORETSE_AHBiiO1I,
output
[
79
:
0
]
CORETSE_AHBOOI1I,
output
CORETSE_AHBol0,
output
CORETSE_AHBil0,
output
CORETSE_AHBO00,
output
CORETSE_AHBI00,
output
CORETSE_AHBIOI1I,
output
[
79
:
0
]
CORETSE_AHBlOI1I,
output
CORETSE_AHBoOI1I
)
;
localparam
CORETSE_AHBiOI1I
=
27
'b
111011100110101100100111110
;
localparam
CORETSE_AHBOII1I
=
28
'b
1110111001101011001001111110
;
reg
[
31
:
0
]
CORETSE_AHBIII1I
;
wire
[
31
:
0
]
CORETSE_AHBlII1I
;
reg
[
47
:
0
]
CORETSE_AHBoII1I
;
wire
[
47
:
0
]
CORETSE_AHBiII1I
;
reg
[
79
:
0
]
CORETSE_AHBOlI1I
;
wire
[
79
:
0
]
CORETSE_AHBIlI1I
;
reg
[
79
:
0
]
CORETSE_AHBllI1I
;
wire
[
79
:
0
]
CORETSE_AHBolI1I
;
reg
CORETSE_AHBilI1I
;
reg
CORETSE_AHBO0I1I
;
reg
CORETSE_AHBI0I1I
;
reg
CORETSE_AHBl0I1I
;
reg
CORETSE_AHBo0I1I
;
reg
CORETSE_AHBi0I1I
;
reg
CORETSE_AHBO1I1I
;
reg
CORETSE_AHBI1I1I
;
reg
CORETSE_AHBl1I1I
;
reg
CORETSE_AHBo1I1I
;
reg
CORETSE_AHBi1I1I
;
reg
CORETSE_AHBOoI1I
;
reg
CORETSE_AHBIoI1I
;
reg
CORETSE_AHBloI1I
;
reg
CORETSE_AHBooI1I
;
wire
CORETSE_AHBioI1I
;
reg
CORETSE_AHBOiI1I
;
wire
CORETSE_AHBIiI1I
;
wire
CORETSE_AHBliI1I
;
wire
CORETSE_AHBoiI1I
;
wire
[
79
:
0
]
CORETSE_AHBiiI1I
;
reg
CORETSE_AHBOOl1I
;
wire
CORETSE_AHBIOl1I
;
wire
CORETSE_AHBlOl1I
;
wire
CORETSE_AHBoOl1I
;
wire
CORETSE_AHBiOl1I
;
reg
CORETSE_AHBOIl1I
;
wire
CORETSE_AHBIIl1I
;
reg
[
7
:
0
]
CORETSE_AHBlIl1I
;
wire
[
7
:
0
]
CORETSE_AHBoIl1I
;
wire
CORETSE_AHBiIl1I
;
reg
CORETSE_AHBOll1I
;
wire
CORETSE_AHBIll1I
;
reg
[
7
:
0
]
CORETSE_AHBlll1I
;
wire
[
7
:
0
]
CORETSE_AHBoll1I
;
wire
CORETSE_AHBill1I
;
reg
CORETSE_AHBO0l1I
;
wire
CORETSE_AHBI0l1I
;
reg
CORETSE_AHBl0l1I
;
wire
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
CORETSE_AHBo0l1I
;
wire
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
CORETSE_AHBi0l1I
;
wire
CORETSE_AHBO1l1I
;
reg
CORETSE_AHBI1l1I
;
reg
CORETSE_AHBl1l1I
;
reg
CORETSE_AHBo1l1I
;
wire
CORETSE_AHBi1l1I
;
wire
[
79
:
0
]
CORETSE_AHBOol1I
;
wire
CORETSE_AHBIol1I
;
reg
CORETSE_AHBlol1I
;
reg
CORETSE_AHBool1I
;
wire
CORETSE_AHBiol1I
;
wire
CORETSE_AHBOil1I
;
wire
CORETSE_AHBIil1I
;
wire
CORETSE_AHBlil1I
;
wire
[
`CORETSE_AHBi1I0
:
`CORETSE_AHBo1I0
]
CORETSE_AHBoil1I
;
wire
[
`CORETSE_AHBIoI0
:
`CORETSE_AHBOoI0
]
CORETSE_AHBiil1I
;
reg
[
23
:
0
]
CORETSE_AHBOO01I
;
wire
[
23
:
0
]
CORETSE_AHBIO01I
;
assign
CORETSE_AHBlil1I
=
CORETSE_AHBOiO1I
[
`CORETSE_AHBl1I0
]
;
assign
CORETSE_AHBoil1I
=
CORETSE_AHBOiO1I
[
`CORETSE_AHBi1I0
:
`CORETSE_AHBo1I0
]
;
assign
CORETSE_AHBiil1I
=
CORETSE_AHBOiO1I
[
`CORETSE_AHBIoI0
:
`CORETSE_AHBOoI0
]
;
assign
CORETSE_AHBoiO1I
=
CORETSE_AHBOiI1I
;
assign
CORETSE_AHBiiO1I
=
CORETSE_AHBOlI1I
;
assign
CORETSE_AHBOOI1I
=
CORETSE_AHBllI1I
;
assign
CORETSE_AHBoOl1I
=
CORETSE_AHBoOo0I
&
CORETSE_AHBi0O1I
;
assign
CORETSE_AHBll0
=
CORETSE_AHBooI1I
;
assign
CORETSE_AHBO00
=
CORETSE_AHBO0l1I
;
assign
CORETSE_AHBI00
=
CORETSE_AHBl0l1I
;
assign
CORETSE_AHBIOI1I
=
CORETSE_AHBi1l1I
;
assign
CORETSE_AHBoOI1I
=
CORETSE_AHBI1l1I
;
assign
CORETSE_AHBiol1I
=
(
~
CORETSE_AHBl0I
&
CORETSE_AHBlol1I
)
|
(
CORETSE_AHBl0I
&
CORETSE_AHBOil1I
)
;
assign
CORETSE_AHBliO1I
=
CORETSE_AHBiol1I
;
assign
CORETSE_AHBOil1I
=
CORETSE_AHBOo0lI
|
CORETSE_AHBlOo0I
;
assign
CORETSE_AHBi1l1I
=
CORETSE_AHBI1I1I
&
(
~
CORETSE_AHBl1I1I
)
;
assign
CORETSE_AHBOol1I
=
{
80
{
CORETSE_AHBO1O1I
&
~
CORETSE_AHBIiO1I
}
}
&
(
CORETSE_AHBI1O1I
+
80
'h
8
)
|
{
80
{
CORETSE_AHBO1O1I
&
CORETSE_AHBIiO1I
}
}
&
(
CORETSE_AHBI1O1I
)
|
{
80
{
~
CORETSE_AHBO1O1I
&
~
CORETSE_AHBIiO1I
}
}
&
(
CORETSE_AHBI1O1I
+
80
'h
10
)
|
{
80
{
~
CORETSE_AHBO1O1I
&
CORETSE_AHBIiO1I
}
}
&
(
CORETSE_AHBI1O1I
)
;
assign
CORETSE_AHBIol1I
=
CORETSE_AHBi1I1I
&
~
CORETSE_AHBOoI1I
;
assign
CORETSE_AHBlOl1I
=
~
CORETSE_AHBIiO1I
&
(
~
CORETSE_AHBioO1I
&
CORETSE_AHBi1l1I
&
CORETSE_AHBi1I1I
&
CORETSE_AHBloI1I
|
CORETSE_AHBioO1I
&
CORETSE_AHBIol1I
&
CORETSE_AHBloI1I
)
|
CORETSE_AHBIiO1I
&
(
CORETSE_AHBOoI1I
&
CORETSE_AHBOOl1I
)
;
assign
CORETSE_AHBIiI1I
=
CORETSE_AHBlOl1I
|
~
CORETSE_AHBlOl1I
&
CORETSE_AHBi1I1I
&
CORETSE_AHBOiI1I
;
assign
CORETSE_AHBiiI1I
=
{
CORETSE_AHBoII1I
,
CORETSE_AHBIII1I
}
;
assign
CORETSE_AHBliI1I
=
CORETSE_AHBO0I1I
&
~
CORETSE_AHBI0I1I
;
assign
CORETSE_AHBoiI1I
=
CORETSE_AHBo0I1I
&
~
CORETSE_AHBi0I1I
;
assign
CORETSE_AHBlOI1I
=
CORETSE_AHBiiI1I
;
assign
CORETSE_AHBIO01I
=
{
24
{
CORETSE_AHBlil1I
}
}
&
(
{
24
{
(
CORETSE_AHBOO01I
==
CORETSE_AHBiil1I
)
}
}
&
24
'b
0
|
{
24
{
!
(
CORETSE_AHBOO01I
==
CORETSE_AHBiil1I
)
}
}
&
(
CORETSE_AHBOO01I
+
1
'b
1
)
)
;
assign
CORETSE_AHBIil1I
=
CORETSE_AHBlil1I
&
(
CORETSE_AHBOO01I
==
CORETSE_AHBiil1I
)
;
assign
CORETSE_AHBlII1I
=
{
32
{
CORETSE_AHBoOl1I
}
}
&
(
{
32
{
(
CORETSE_AHBlOl1I
&
~
CORETSE_AHBIiO1I
)
}
}
&
CORETSE_AHBOol1I
[
31
:
0
]
|
{
32
{
(
CORETSE_AHBlOl1I
&
CORETSE_AHBIiO1I
&
~
CORETSE_AHBO1O1I
)
}
}
&
(
CORETSE_AHBOol1I
[
31
:
0
]
+
{
29
'b
0
,
CORETSE_AHBIII1I
[
2
:
0
]
}
)
|
{
32
{
(
CORETSE_AHBlOl1I
&
CORETSE_AHBIiO1I
&
CORETSE_AHBO1O1I
)
}
}
&
(
CORETSE_AHBOol1I
[
31
:
0
]
+
{
30
'b
0
,
CORETSE_AHBIII1I
[
1
:
0
]
}
)
|
{
32
{
(
~
CORETSE_AHBlOl1I
&
CORETSE_AHBIil1I
&
~
CORETSE_AHBOOl1I
)
}
}
&
(
{
24
'b
0
,
CORETSE_AHBoil1I
}
+
CORETSE_AHBIII1I
[
31
:
0
]
)
|
{
32
{
(
~
CORETSE_AHBlOl1I
&
CORETSE_AHBIil1I
&
CORETSE_AHBOOl1I
)
}
}
&
{
24
'b
0
,
CORETSE_AHBoil1I
}
|
{
32
{
(
~
CORETSE_AHBlOl1I
&
~
CORETSE_AHBIil1I
&
CORETSE_AHBOOl1I
&
~
CORETSE_AHBO1O1I
)
}
}
&
{
29
'b
0
,
CORETSE_AHBIII1I
[
2
:
0
]
}
|
{
32
{
(
~
CORETSE_AHBlOl1I
&
~
CORETSE_AHBIil1I
&
CORETSE_AHBOOl1I
&
CORETSE_AHBO1O1I
)
}
}
&
{
30
'b
0
,
CORETSE_AHBIII1I
[
1
:
0
]
}
|
{
32
{
(
~
CORETSE_AHBlOl1I
&
~
CORETSE_AHBIil1I
&
~
CORETSE_AHBOOl1I
&
~
CORETSE_AHBO1O1I
)
}
}
&
(
CORETSE_AHBIII1I
+
32
'h
8
)
|
{
32
{
(
~
CORETSE_AHBlOl1I
&
~
CORETSE_AHBIil1I
&
~
CORETSE_AHBOOl1I
&
CORETSE_AHBO1O1I
)
}
}
&
(
CORETSE_AHBIII1I
+
32
'h
4
)
)
;
assign
CORETSE_AHBIOl1I
=
~
CORETSE_AHBOOl1I
&
(
~
CORETSE_AHBO1O1I
&
~
CORETSE_AHBIII1I
[
31
]
&
(
CORETSE_AHBIII1I
[
29
:
3
]
>=
CORETSE_AHBiOI1I
)
|
CORETSE_AHBO1O1I
&
~
CORETSE_AHBIII1I
[
31
]
&
(
CORETSE_AHBIII1I
[
29
:
2
]
>=
CORETSE_AHBOII1I
)
)
;
assign
CORETSE_AHBiII1I
=
{
48
{
CORETSE_AHBoOl1I
}
}
&
(
(
{
48
{
CORETSE_AHBlOl1I
&
~
CORETSE_AHBIiO1I
}
}
&
CORETSE_AHBOol1I
[
79
:
32
]
)
|
(
{
48
{
CORETSE_AHBlOl1I
&
CORETSE_AHBIiO1I
}
}
&
(
CORETSE_AHBoII1I
+
CORETSE_AHBOol1I
[
79
:
32
]
+
1
'b
1
)
)
|
(
{
48
{
~
CORETSE_AHBlOl1I
&
CORETSE_AHBOOl1I
}
}
&
(
CORETSE_AHBoII1I
+
1
'b
1
)
)
|
(
{
48
{
~
CORETSE_AHBlOl1I
&
~
CORETSE_AHBOOl1I
}
}
&
CORETSE_AHBoII1I
)
)
;
assign
CORETSE_AHBioI1I
=
~
CORETSE_AHBOOl1I
&
CORETSE_AHBooI1I
|
CORETSE_AHBOOl1I
&
~
CORETSE_AHBooI1I
;
assign
CORETSE_AHBO1l1I
=
CORETSE_AHBl1l1I
&
1
'b
0
|
~
CORETSE_AHBl1l1I
&
CORETSE_AHBOOl1I
&
1
'b
1
|
~
CORETSE_AHBl1l1I
&
~
CORETSE_AHBOOl1I
&
CORETSE_AHBI1l1I
;
assign
CORETSE_AHBIlI1I
=
(
{
80
{
CORETSE_AHBliI1I
}
}
&
CORETSE_AHBiiI1I
)
|
(
{
80
{
~
CORETSE_AHBliI1I
}
}
&
CORETSE_AHBOlI1I
)
;
assign
CORETSE_AHBolI1I
=
(
{
80
{
CORETSE_AHBoiI1I
}
}
&
CORETSE_AHBiiI1I
)
|
(
{
80
{
~
CORETSE_AHBoiI1I
}
}
&
CORETSE_AHBllI1I
)
;
assign
CORETSE_AHBiOl1I
=
CORETSE_AHBO1O1I
&
CORETSE_AHBO0O1I
&
(
CORETSE_AHBl0O1I
[
79
:
2
]
==
CORETSE_AHBiiI1I
[
79
:
2
]
)
|
~
CORETSE_AHBO1O1I
&
CORETSE_AHBO0O1I
&
(
CORETSE_AHBl0O1I
[
79
:
3
]
==
CORETSE_AHBiiI1I
[
79
:
3
]
)
;
assign
CORETSE_AHBoIl1I
=
{
8
{
CORETSE_AHBiOl1I
&
~
CORETSE_AHBOIl1I
}
}
&
8
'b
00000001
|
{
8
{
CORETSE_AHBOIl1I
}
}
&
(
CORETSE_AHBlIl1I
+
1
'b
1
)
|
{
8
{
~
CORETSE_AHBiOl1I
&
~
CORETSE_AHBOIl1I
}
}
&
CORETSE_AHBlIl1I
;
assign
CORETSE_AHBIIl1I
=
CORETSE_AHBiOl1I
&
1
'b
1
|
~
CORETSE_AHBiOl1I
&
(
CORETSE_AHBlIl1I
==
CORETSE_AHBolO1I
)
&
1
'b
0
|
~
CORETSE_AHBiOl1I
&
~
(
CORETSE_AHBlIl1I
==
CORETSE_AHBolO1I
)
&
CORETSE_AHBOIl1I
;
assign
CORETSE_AHBol0
=
CORETSE_AHBOIl1I
;
assign
CORETSE_AHBiIl1I
=
CORETSE_AHBO1O1I
&
CORETSE_AHBI0O1I
&
(
CORETSE_AHBo0O1I
[
79
:
2
]
==
CORETSE_AHBiiI1I
[
79
:
2
]
)
|
~
CORETSE_AHBO1O1I
&
CORETSE_AHBI0O1I
&
(
CORETSE_AHBo0O1I
[
79
:
3
]
==
CORETSE_AHBiiI1I
[
79
:
3
]
)
;
assign
CORETSE_AHBoll1I
=
{
8
{
CORETSE_AHBiIl1I
&
~
CORETSE_AHBOll1I
}
}
&
8
'b
00000001
|
{
8
{
CORETSE_AHBOll1I
}
}
&
(
CORETSE_AHBlll1I
+
1
'b
1
)
|
{
8
{
~
CORETSE_AHBiIl1I
&
~
CORETSE_AHBOll1I
}
}
&
CORETSE_AHBlll1I
;
assign
CORETSE_AHBIll1I
=
CORETSE_AHBiIl1I
&
1
'b
1
|
~
CORETSE_AHBiIl1I
&
(
CORETSE_AHBlll1I
==
CORETSE_AHBilO1I
)
&
1
'b
0
|
~
CORETSE_AHBiIl1I
&
~
(
CORETSE_AHBlll1I
==
CORETSE_AHBilO1I
)
&
CORETSE_AHBOll1I
;
assign
CORETSE_AHBil0
=
CORETSE_AHBOll1I
;
genvar
CORETSE_AHBOloI
;
generate
for
(
CORETSE_AHBOloI
=
0
;
CORETSE_AHBOloI
<=
(
CORETSE_AHBlII
-
CORETSE_AHBIII
)
;
CORETSE_AHBOloI
=
CORETSE_AHBOloI
+
1
)
begin
:
CORETSE_AHBlO01I
assign
CORETSE_AHBo0l1I
[
CORETSE_AHBOloI
]
=
~
CORETSE_AHBO1O1I
&
CORETSE_AHBiiI1I
[
CORETSE_AHBIII
+
2
+
CORETSE_AHBOloI
]
&
CORETSE_AHBloO1I
[
CORETSE_AHBOloI
]
|
CORETSE_AHBO1O1I
&
CORETSE_AHBiiI1I
[
CORETSE_AHBIII
+
1
+
CORETSE_AHBOloI
]
&
CORETSE_AHBloO1I
[
CORETSE_AHBOloI
]
;
end
assign
CORETSE_AHBill1I
=
|
CORETSE_AHBo0l1I
;
endgenerate
genvar
CORETSE_AHBoO01I
;
generate
for
(
CORETSE_AHBoO01I
=
0
;
CORETSE_AHBoO01I
<=
(
CORETSE_AHBiII
-
CORETSE_AHBoII
)
;
CORETSE_AHBoO01I
=
CORETSE_AHBoO01I
+
1
)
begin
:
CORETSE_AHBiO01I
assign
CORETSE_AHBi0l1I
[
CORETSE_AHBoO01I
]
=
~
CORETSE_AHBO1O1I
&
CORETSE_AHBiiI1I
[
CORETSE_AHBoII
+
2
+
CORETSE_AHBoO01I
]
&
CORETSE_AHBooO1I
[
CORETSE_AHBoO01I
]
|
CORETSE_AHBO1O1I
&
CORETSE_AHBiiI1I
[
CORETSE_AHBoII
+
1
+
CORETSE_AHBoO01I
]
&
CORETSE_AHBooO1I
[
CORETSE_AHBoO01I
]
;
end
assign
CORETSE_AHBI0l1I
=
|
CORETSE_AHBi0l1I
;
endgenerate
always
@
(
posedge
CORETSE_AHBOl0
or
posedge
CORETSE_AHBiol1I
)
begin
if
(
CORETSE_AHBiol1I
)
begin
CORETSE_AHBilI1I
<=
1
'b
0
;
CORETSE_AHBO0I1I
<=
1
'b
0
;
CORETSE_AHBI0I1I
<=
1
'b
0
;
CORETSE_AHBl0I1I
<=
1
'b
0
;
CORETSE_AHBo0I1I
<=
1
'b
0
;
CORETSE_AHBi0I1I
<=
1
'b
0
;
CORETSE_AHBO1I1I
<=
1
'b
0
;
CORETSE_AHBI1I1I
<=
1
'b
0
;
CORETSE_AHBl1I1I
<=
1
'b
0
;
CORETSE_AHBo1I1I
<=
1
'b
0
;
CORETSE_AHBi1I1I
<=
1
'b
0
;
CORETSE_AHBOoI1I
<=
1
'b
0
;
CORETSE_AHBIoI1I
<=
1
'b
0
;
CORETSE_AHBloI1I
<=
1
'b
0
;
CORETSE_AHBo1l1I
<=
1
'b
0
;
CORETSE_AHBl1l1I
<=
1
'b
0
;
CORETSE_AHBOlI1I
<=
80
'b
0
;
CORETSE_AHBllI1I
<=
80
'b
0
;
CORETSE_AHBoII1I
<=
48
'b
0
;
CORETSE_AHBIII1I
<=
32
'b
0
;
CORETSE_AHBOiI1I
<=
1
'b
0
;
CORETSE_AHBI1l1I
<=
1
'b
0
;
CORETSE_AHBooI1I
<=
1
'b
0
;
CORETSE_AHBOIl1I
<=
1
'b
0
;
CORETSE_AHBOll1I
<=
1
'b
0
;
CORETSE_AHBlIl1I
<=
8
'b
0
;
CORETSE_AHBlll1I
<=
8
'b
0
;
CORETSE_AHBO0l1I
<=
1
'b
0
;
CORETSE_AHBl0l1I
<=
1
'b
0
;
CORETSE_AHBOO01I
<=
24
'b
0
;
CORETSE_AHBOOl1I
<=
1
'b
0
;
end
else
begin
CORETSE_AHBilI1I
<=
CORETSE_AHBi1O1I
;
CORETSE_AHBO0I1I
<=
CORETSE_AHBilI1I
;
CORETSE_AHBI0I1I
<=
CORETSE_AHBO0I1I
;
CORETSE_AHBl0I1I
<=
CORETSE_AHBOoO1I
;
CORETSE_AHBo0I1I
<=
CORETSE_AHBl0I1I
;
CORETSE_AHBi0I1I
<=
CORETSE_AHBo0I1I
;
CORETSE_AHBO1I1I
<=
CORETSE_AHBIl0
;
CORETSE_AHBI1I1I
<=
CORETSE_AHBO1I1I
;
CORETSE_AHBl1I1I
<=
CORETSE_AHBI1I1I
;
CORETSE_AHBo1I1I
<=
CORETSE_AHBl1O1I
;
CORETSE_AHBi1I1I
<=
CORETSE_AHBo1I1I
;
CORETSE_AHBOoI1I
<=
CORETSE_AHBi1I1I
;
CORETSE_AHBIoI1I
<=
CORETSE_AHBo1O1I
;
CORETSE_AHBloI1I
<=
CORETSE_AHBIoI1I
;
CORETSE_AHBo1l1I
<=
CORETSE_AHBIoO1I
;
CORETSE_AHBl1l1I
<=
CORETSE_AHBo1l1I
;
CORETSE_AHBOlI1I
<=
CORETSE_AHBIlI1I
;
CORETSE_AHBllI1I
<=
CORETSE_AHBolI1I
;
CORETSE_AHBoII1I
<=
CORETSE_AHBiII1I
;
CORETSE_AHBIII1I
<=
CORETSE_AHBlII1I
;
CORETSE_AHBOiI1I
<=
CORETSE_AHBIiI1I
;
CORETSE_AHBI1l1I
<=
CORETSE_AHBO1l1I
;
CORETSE_AHBooI1I
<=
CORETSE_AHBioI1I
;
CORETSE_AHBOIl1I
<=
CORETSE_AHBIIl1I
;
CORETSE_AHBOll1I
<=
CORETSE_AHBIll1I
;
CORETSE_AHBlIl1I
<=
CORETSE_AHBoIl1I
;
CORETSE_AHBlll1I
<=
CORETSE_AHBoll1I
;
CORETSE_AHBO0l1I
<=
CORETSE_AHBill1I
;
CORETSE_AHBl0l1I
<=
CORETSE_AHBI0l1I
;
CORETSE_AHBOO01I
<=
CORETSE_AHBIO01I
;
CORETSE_AHBOOl1I
<=
CORETSE_AHBIOl1I
;
end
end
always
@
(
posedge
CORETSE_AHBOl0
or
posedge
CORETSE_AHBOil1I
)
begin
if
(
CORETSE_AHBOil1I
)
begin
CORETSE_AHBool1I
<=
1
'b
1
;
CORETSE_AHBlol1I
<=
1
'b
1
;
end
else
begin
CORETSE_AHBool1I
<=
1
'b
0
;
CORETSE_AHBlol1I
<=
CORETSE_AHBool1I
;
end
end
endmodule
