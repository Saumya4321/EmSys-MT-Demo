// VERSION     : $Revision: 1.5 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
petmc_top
(
CORETSE_AHBiOO1
,
CORETSE_AHBo1Oo
,
CORETSE_AHBiio
,
CORETSE_AHBiOi
,
CORETSE_AHBIIi
,
CORETSE_AHBOIi
,
CORETSE_AHBoOi
,
CORETSE_AHBl0Io
,
CORETSE_AHBo0Io
,
CORETSE_AHBi0Io
,
CORETSE_AHBO1Io
,
CORETSE_AHBoIi1
,
CORETSE_AHBoo01
,
CORETSE_AHBll00
,
CORETSE_AHBlIi
,
CORETSE_AHBi111
,
CORETSE_AHBOoOo
,
CORETSE_AHBOiIo
,
CORETSE_AHBo0Oo
,
CORETSE_AHBOlIo
,
CORETSE_AHBIlIo
,
CORETSE_AHBllIo
,
CORETSE_AHBolIo
,
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
,
CORETSE_AHBIoo
,
CORETSE_AHBo0o1
,
CORETSE_AHBoOo1
,
CORETSE_AHBilIo
,
CORETSE_AHBO0Io
)
;
input
CORETSE_AHBiOO1
,
CORETSE_AHBo1Oo
;
input
[
7
:
0
]
CORETSE_AHBiio
;
input
CORETSE_AHBiOi
,
CORETSE_AHBIIi
,
CORETSE_AHBOIi
,
CORETSE_AHBoOi
;
input
CORETSE_AHBl0Io
,
CORETSE_AHBo0Io
,
CORETSE_AHBi0Io
,
CORETSE_AHBO1Io
;
input
CORETSE_AHBoIi1
;
input
[
1
:
0
]
CORETSE_AHBoo01
;
input
[
47
:
0
]
CORETSE_AHBll00
;
input
CORETSE_AHBlIi
;
input
[
15
:
0
]
CORETSE_AHBi111
,
CORETSE_AHBOoOo
;
input
CORETSE_AHBOiIo
;
input
CORETSE_AHBo0Oo
;
output
[
7
:
0
]
CORETSE_AHBOlIo
;
output
CORETSE_AHBIlIo
,
CORETSE_AHBllIo
,
CORETSE_AHBolIo
;
output
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
;
output
CORETSE_AHBIoo
;
output
CORETSE_AHBoOo1
,
CORETSE_AHBilIo
,
CORETSE_AHBO0Io
;
output
[
7
:
0
]
CORETSE_AHBo0o1
;
reg
[
7
:
0
]
CORETSE_AHBOlIo
;
reg
CORETSE_AHBIlIo
,
CORETSE_AHBllIo
,
CORETSE_AHBolIo
;
reg
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
;
reg
CORETSE_AHBIoo
;
reg
CORETSE_AHBoOo1
,
CORETSE_AHBilIo
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBoollI
,
CORETSE_AHBiollI
,
CORETSE_AHBOillI
;
reg
CORETSE_AHBIillI
,
CORETSE_AHBlillI
;
wire
CORETSE_AHBoillI
;
reg
CORETSE_AHBiillI
;
wire
CORETSE_AHBOO0lI
,
CORETSE_AHBIO0lI
,
CORETSE_AHBI1llI
,
CORETSE_AHBlO0lI
;
reg
CORETSE_AHBO0Io
,
CORETSE_AHBoO0lI
,
CORETSE_AHBo1llI
,
CORETSE_AHBiO0lI
;
wire
[
5
:
0
]
CORETSE_AHBOI0lI
;
wire
CORETSE_AHBII0lI
,
CORETSE_AHBlI0lI
;
wire
[
5
:
0
]
CORETSE_AHBoI0lI
;
reg
[
5
:
0
]
CORETSE_AHBiI0lI
;
wire
[
7
:
0
]
CORETSE_AHBOl0lI
;
wire
[
7
:
0
]
CORETSE_AHBIl0lI
;
wire
CORETSE_AHBll0lI
,
CORETSE_AHBol0lI
,
CORETSE_AHBil0lI
;
wire
CORETSE_AHBO00lI
,
CORETSE_AHBI00lI
,
CORETSE_AHBl00lI
;
reg
CORETSE_AHBo00lI
,
CORETSE_AHBi00lI
,
CORETSE_AHBO10lI
;
wire
CORETSE_AHBliOlI
,
CORETSE_AHBoiOlI
,
CORETSE_AHBiiOlI
,
CORETSE_AHBOOIlI
;
wire
CORETSE_AHBI10lI
;
wire
CORETSE_AHBl10lI
,
CORETSE_AHBo10lI
;
assign
CORETSE_AHBo0o1
=
CORETSE_AHBIl0lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBoollI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoollI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIi1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBiollI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiollI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoollI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBOillI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOillI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiollI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBIillI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIillI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiIo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBlillI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBlillI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIillI
;
end
assign
CORETSE_AHBoillI
=
~
CORETSE_AHBiillI
&
CORETSE_AHBlIi
&
CORETSE_AHBoIi1
&
CORETSE_AHBIoo
|
CORETSE_AHBiillI
&
~
(
CORETSE_AHBiO0lI
&
CORETSE_AHBo0Io
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBiillI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiillI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoillI
;
end
assign
CORETSE_AHBOO0lI
=
CORETSE_AHBoO0lI
&
CORETSE_AHBI1llI
&
~
CORETSE_AHBo1llI
|
CORETSE_AHBO0Io
&
~
(
CORETSE_AHBiOi
&
(
~
CORETSE_AHBlillI
|
CORETSE_AHBoOi
)
|
CORETSE_AHBiillI
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBO0Io
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO0Io
<=
#
CORETSE_AHBIoII
CORETSE_AHBOO0lI
;
end
assign
CORETSE_AHBIO0lI
=
CORETSE_AHBO0Io
&
(
CORETSE_AHBiOi
&
(
~
CORETSE_AHBlillI
|
CORETSE_AHBoOi
)
|
CORETSE_AHBiillI
)
|
CORETSE_AHBoO0lI
&
~
(
CORETSE_AHBI1llI
&
~
CORETSE_AHBo1llI
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBoO0lI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoO0lI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIO0lI
;
end
assign
CORETSE_AHBI1llI
=
~
CORETSE_AHBiO0lI
&
(
CORETSE_AHBOOo1
|
CORETSE_AHBilo
)
|
CORETSE_AHBiO0lI
&
CORETSE_AHBo0Io
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBo1llI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBo1llI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1llI
;
end
assign
CORETSE_AHBlO0lI
=
CORETSE_AHBO0Io
&
CORETSE_AHBiillI
|
CORETSE_AHBoO0lI
&
CORETSE_AHBiO0lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBiO0lI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiO0lI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO0lI
;
end
assign
CORETSE_AHBII0lI
=
~
CORETSE_AHBiO0lI
|
CORETSE_AHBiO0lI
&
CORETSE_AHBiI0lI
[
5
:
0
]
==
6
'h
13
&
(
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBi00lI
|
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBO10lI
)
;
assign
CORETSE_AHBOI0lI
[
5
:
0
]
=
6
'h
00
;
assign
CORETSE_AHBlI0lI
=
CORETSE_AHBiO0lI
&
CORETSE_AHBiI0lI
[
5
:
0
]
!=
6
'h
14
&
(
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBi00lI
|
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBO10lI
)
;
assign
CORETSE_AHBoI0lI
[
5
:
0
]
=
{
6
{
CORETSE_AHBII0lI
}
}
&
CORETSE_AHBOI0lI
[
5
:
0
]
|
{
6
{
~
CORETSE_AHBII0lI
&
CORETSE_AHBlI0lI
}
}
&
CORETSE_AHBiI0lI
[
5
:
0
]
+
1
'b
1
|
{
6
{
~
CORETSE_AHBII0lI
&
~
CORETSE_AHBlI0lI
}
}
&
CORETSE_AHBiI0lI
[
5
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBiI0lI
[
5
:
0
]
<=
#
CORETSE_AHBIoII
6
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiI0lI
[
5
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI0lI
[
5
:
0
]
;
end
assign
CORETSE_AHBOl0lI
[
7
:
0
]
=
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
00
}
}
&
8
'h
01
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
01
}
}
&
8
'h
80
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
02
}
}
&
8
'h
c2
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
03
}
}
&
8
'h
00
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
04
}
}
&
8
'h
00
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
05
}
}
&
8
'h
01
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
06
}
}
&
CORETSE_AHBll00
[
47
:
40
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
07
}
}
&
CORETSE_AHBll00
[
39
:
32
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
08
}
}
&
CORETSE_AHBll00
[
31
:
24
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
09
}
}
&
CORETSE_AHBll00
[
23
:
16
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
0a
}
}
&
CORETSE_AHBll00
[
15
:
8
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
0b
}
}
&
CORETSE_AHBll00
[
7
:
0
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
0c
}
}
&
8
'h
88
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
0d
}
}
&
8
'h
08
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
0e
}
}
&
8
'h
00
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
0f
}
}
&
8
'h
01
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
10
}
}
&
CORETSE_AHBi111
[
15
:
8
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
11
}
}
&
CORETSE_AHBi111
[
7
:
0
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
12
}
}
&
CORETSE_AHBOoOo
[
15
:
8
]
|
{
8
{
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
13
}
}
&
CORETSE_AHBOoOo
[
7
:
0
]
;
assign
CORETSE_AHBIl0lI
[
7
:
0
]
=
{
8
{
~
CORETSE_AHBiO0lI
}
}
&
CORETSE_AHBiio
[
7
:
0
]
|
{
8
{
CORETSE_AHBiO0lI
}
}
&
CORETSE_AHBOl0lI
[
7
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBOlIo
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOlIo
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl0lI
[
7
:
0
]
;
end
assign
CORETSE_AHBll0lI
=
~
CORETSE_AHBiO0lI
&
CORETSE_AHBoO0lI
&
CORETSE_AHBiOi
|
CORETSE_AHBiO0lI
&
CORETSE_AHBoO0lI
&
CORETSE_AHBiillI
|
CORETSE_AHBiO0lI
&
CORETSE_AHBIlIo
&
~
CORETSE_AHBi00lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBIlIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIlIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBll0lI
;
end
assign
CORETSE_AHBO00lI
=
CORETSE_AHBiO0lI
&
CORETSE_AHBl0Io
&
~
CORETSE_AHBOIi
&
~
CORETSE_AHBolIo
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBo00lI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBo00lI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO00lI
;
end
assign
CORETSE_AHBI00lI
=
CORETSE_AHBo00lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBi00lI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi00lI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI00lI
;
end
assign
CORETSE_AHBl00lI
=
CORETSE_AHBi00lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBO10lI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO10lI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00lI
;
end
assign
CORETSE_AHBol0lI
=
~
CORETSE_AHBiO0lI
&
CORETSE_AHBIIi
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBllIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBllIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0lI
;
end
assign
CORETSE_AHBil0lI
=
~
CORETSE_AHBiO0lI
&
CORETSE_AHBOIi
|
CORETSE_AHBiO0lI
&
CORETSE_AHBiI0lI
[
4
:
0
]
==
5
'h
13
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBolIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBolIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBil0lI
;
end
assign
CORETSE_AHBliOlI
=
~
CORETSE_AHBiO0lI
&
CORETSE_AHBl0Io
&
~
CORETSE_AHBOIi
&
~
CORETSE_AHBolIo
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBolo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBolo
<=
#
CORETSE_AHBIoII
CORETSE_AHBliOlI
;
end
assign
CORETSE_AHBoiOlI
=
CORETSE_AHBo0Io
|
CORETSE_AHBiO0lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBOOo1
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiOlI
;
end
assign
CORETSE_AHBiiOlI
=
CORETSE_AHBi0Io
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBO0o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiOlI
;
end
assign
CORETSE_AHBOOIlI
=
CORETSE_AHBO1Io
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBilo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBilo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOIlI
;
end
assign
CORETSE_AHBI10lI
=
~
CORETSE_AHBIoo
&
(
~
CORETSE_AHBl10lI
&
CORETSE_AHBilIo
|
CORETSE_AHBiollI
&
~
CORETSE_AHBOillI
)
|
CORETSE_AHBIoo
&
CORETSE_AHBiollI
&
~
CORETSE_AHBlIi
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBIoo
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIoo
<=
#
CORETSE_AHBIoII
CORETSE_AHBI10lI
;
end
assign
CORETSE_AHBl10lI
=
CORETSE_AHBiO0lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBoOo1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBl10lI
;
end
assign
CORETSE_AHBo10lI
=
CORETSE_AHBiO0lI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBo0Oo
)
begin
if
(
CORETSE_AHBo0Oo
)
CORETSE_AHBilIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBilIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBo10lI
;
end
endmodule
