// REVISION    : $Revision: 1.4 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxtfif_fab
#
(
parameter
TABITS
=
12
,
parameter
CORETSE_AHBIo1
=
32
,
parameter
CORETSE_AHBlo1
=
$clog2
(
CORETSE_AHBIo1
/
8
)
)
(
CORETSE_AHBOOo
,
CORETSE_AHBilII
,
CORETSE_AHBiiOI
,
CORETSE_AHBIOo
,
CORETSE_AHBlOo
,
CORETSE_AHBoOo
,
CORETSE_AHBiOo
,
CORETSE_AHBOIo
,
CORETSE_AHBIIo
,
CORETSE_AHBlIo
,
CORETSE_AHBoIo
,
CORETSE_AHBiIo
,
CORETSE_AHBl1i
,
CORETSE_AHBo1i
,
CORETSE_AHBi1i
,
CORETSE_AHBl1OI
,
CORETSE_AHBo1OI
,
CORETSE_AHBiOII
,
CORETSE_AHBOIII
,
CORETSE_AHBIIII
,
CORETSE_AHBoOOI
,
CORETSE_AHBIli
,
CORETSE_AHBlli
,
CORETSE_AHBOli
,
CORETSE_AHBloo
,
CORETSE_AHBooo
,
CORETSE_AHBOoi
,
CORETSE_AHBIoi
,
CORETSE_AHBloi
,
CORETSE_AHBiIOI
,
CORETSE_AHBOlOI
)
;
input
CORETSE_AHBOOo
;
input
CORETSE_AHBilII
;
input
CORETSE_AHBiiOI
;
input
[
(
CORETSE_AHBIo1
-
1
)
:
0
]
CORETSE_AHBIOo
;
input
CORETSE_AHBlOo
;
input
CORETSE_AHBoOo
;
input
[
1
:
0
]
CORETSE_AHBiOo
;
input
CORETSE_AHBOIo
;
input
CORETSE_AHBIIo
;
input
[
1
:
0
]
CORETSE_AHBlIo
;
input
CORETSE_AHBoIo
;
input
CORETSE_AHBiIo
;
input
CORETSE_AHBl1i
;
input
[
TABITS
:
0
]
CORETSE_AHBo1i
;
input
CORETSE_AHBi1i
;
input
[
TABITS
:
0
]
CORETSE_AHBl1OI
;
input
[
TABITS
:
0
]
CORETSE_AHBo1OI
;
input
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBiOII
;
input
CORETSE_AHBOIII
;
input
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIIII
;
output
CORETSE_AHBoOOI
;
output
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBIli
;
output
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBlli
;
output
CORETSE_AHBOli
;
output
CORETSE_AHBloo
;
output
CORETSE_AHBooo
;
output
[
TABITS
:
0
]
CORETSE_AHBOoi
;
output
CORETSE_AHBIoi
;
output
CORETSE_AHBloi
;
output
CORETSE_AHBiIOI
;
output
[
TABITS
:
0
]
CORETSE_AHBOlOI
;
parameter
CORETSE_AHBoloI
=
{
TABITS
{
1
'b
0
}
}
;
parameter
CORETSE_AHBol0I
=
{
(
TABITS
+
1
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBIoII
=
1
;
reg
[
TABITS
:
0
]
CORETSE_AHBOoi
;
reg
[
TABITS
:
0
]
CORETSE_AHBiloI
;
reg
[
TABITS
:
0
]
CORETSE_AHBO0oI
;
reg
CORETSE_AHBI0oI
;
reg
CORETSE_AHBIoi
;
reg
CORETSE_AHBloi
;
reg
CORETSE_AHBoOOI
;
wire
CORETSE_AHBloo
;
reg
CORETSE_AHBooo
;
wire
CORETSE_AHBO01I
;
wire
CORETSE_AHBl0oI
;
reg
[
TABITS
:
0
]
CORETSE_AHBo0oI
;
reg
CORETSE_AHBi0oI
;
reg
CORETSE_AHBO1oI
;
reg
CORETSE_AHBI1oI
;
reg
CORETSE_AHBl1oI
;
reg
CORETSE_AHBo1oI
;
reg
CORETSE_AHBi1oI
;
reg
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBIli
;
reg
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBlli
;
reg
CORETSE_AHBOli
;
reg
CORETSE_AHBOooI
;
reg
CORETSE_AHBIooI
;
wire
[
TABITS
:
0
]
CORETSE_AHBlooI
;
reg
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBoooI
;
reg
[
TABITS
:
0
]
CORETSE_AHBiooI
;
reg
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBOioI
;
reg
[
TABITS
:
0
]
CORETSE_AHBIioI
;
reg
CORETSE_AHBO10I
;
reg
[
TABITS
:
0
]
CORETSE_AHBlioI
;
reg
CORETSE_AHBoioI
;
wire
[
TABITS
:
0
]
CORETSE_AHBiioI
;
reg
CORETSE_AHBOOiI
;
reg
CORETSE_AHBIOiI
;
wire
CORETSE_AHBlOiI
;
reg
CORETSE_AHBiIOI
;
wire
[
TABITS
:
0
]
CORETSE_AHBOlOI
;
reg
CORETSE_AHBoOiI
;
//      generated as part of synthesis results.
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBIli
<=
#
1000
CORETSE_AHBoloI
;
else
CORETSE_AHBIli
<=
#
1000
(
{
TABITS
{
~
(
~
CORETSE_AHBiOII
[
TABITS
+
1
]
&
CORETSE_AHBlOiI
)
}
}
&
CORETSE_AHBO0oI
[
(
TABITS
-
1
)
:
0
]
)
|
(
{
TABITS
{
(
~
CORETSE_AHBiOII
[
TABITS
+
1
]
&
CORETSE_AHBlOiI
)
}
}
&
CORETSE_AHBiOII
[
(
TABITS
-
1
)
:
0
]
)
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBlli
<=
#
1000
{
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
{
1
'h
0
}
}
;
else
CORETSE_AHBlli
<=
#
1000
(
{
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
{
~
CORETSE_AHBilII
&
~
(
~
CORETSE_AHBiOII
[
TABITS
+
1
]
&
CORETSE_AHBlOiI
)
}
}
&
{
CORETSE_AHBoIo
,
CORETSE_AHBlIo
,
CORETSE_AHBIIo
,
CORETSE_AHBOIo
,
CORETSE_AHBoOo
,
CORETSE_AHBiOo
,
CORETSE_AHBIOo
}
)
|
(
{
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
{
~
CORETSE_AHBilII
&
(
~
CORETSE_AHBiOII
[
TABITS
+
1
]
&
CORETSE_AHBlOiI
)
}
}
&
CORETSE_AHBIIII
)
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBOli
<=
#
1000
1
'b
0
;
else
CORETSE_AHBOli
<=
#
1000
~
(
CORETSE_AHBl0oI
|
(
~
CORETSE_AHBiOII
[
TABITS
+
1
]
&
CORETSE_AHBlOiI
)
)
;
end
assign
CORETSE_AHBO01I
=
(
CORETSE_AHBO0oI
[
(
TABITS
-
1
)
:
0
]
==
CORETSE_AHBo0oI
[
(
TABITS
-
1
)
:
0
]
)
&
(
CORETSE_AHBO0oI
[
TABITS
]
!=
CORETSE_AHBo0oI
[
TABITS
]
)
;
assign
CORETSE_AHBloo
=
~
CORETSE_AHBO01I
&
CORETSE_AHBoOOI
;
assign
CORETSE_AHBl0oI
=
(
CORETSE_AHBiIo
&
CORETSE_AHBloo
)
;
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBO0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBiOII
[
TABITS
+
1
]
&
CORETSE_AHBlOiI
)
CORETSE_AHBO0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOII
[
TABITS
:
0
]
;
else
if
(
CORETSE_AHBl0oI
)
CORETSE_AHBO0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
+
1
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBo0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBl1oI
&
~
CORETSE_AHBloi
)
CORETSE_AHBo0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1i
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBOooI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
[
TABITS
]
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBIooI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0oI
[
TABITS
]
;
end
assign
CORETSE_AHBlooI
=
(
CORETSE_AHBOooI
==
CORETSE_AHBIooI
)
?
{
1
'b
0
,
CORETSE_AHBoooI
}
:
CORETSE_AHBiooI
;
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBooo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBooo
<=
#
CORETSE_AHBIoII
(
CORETSE_AHBlooI
>
CORETSE_AHBl1OI
)
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBoooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoloI
;
else
CORETSE_AHBoooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
[
(
TABITS
-
1
)
:
0
]
-
CORETSE_AHBo0oI
[
(
TABITS
-
1
)
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBiooI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
CORETSE_AHBiooI
<=
#
CORETSE_AHBIoII
{
1
'b
1
,
CORETSE_AHBO0oI
[
(
TABITS
-
1
)
:
0
]
}
-
{
1
'b
0
,
CORETSE_AHBo0oI
[
(
TABITS
-
1
)
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBlioI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBoOo
&
CORETSE_AHBl0oI
)
CORETSE_AHBlioI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBOioI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoloI
;
else
CORETSE_AHBOioI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
[
(
TABITS
-
1
)
:
0
]
-
CORETSE_AHBlioI
[
(
TABITS
-
1
)
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBIioI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
CORETSE_AHBIioI
<=
#
CORETSE_AHBIoII
{
1
'b
1
,
CORETSE_AHBO0oI
[
(
TABITS
-
1
)
:
0
]
}
-
{
1
'b
0
,
CORETSE_AHBlioI
[
(
TABITS
-
1
)
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBoioI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoioI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlioI
[
TABITS
]
;
end
assign
CORETSE_AHBiioI
=
(
CORETSE_AHBOooI
==
CORETSE_AHBoioI
)
?
{
1
'b
0
,
CORETSE_AHBOioI
}
:
CORETSE_AHBIioI
;
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBoOiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0oI
&
CORETSE_AHBoOo
)
CORETSE_AHBoOiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
(
CORETSE_AHBiioI
>
CORETSE_AHBo1OI
)
&
CORETSE_AHBO10I
)
CORETSE_AHBoOiI
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBiloI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBl0oI
&
(
CORETSE_AHBoOo
|
CORETSE_AHBoOiI
)
)
CORETSE_AHBiloI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
+
1
;
else
if
(
~
CORETSE_AHBO10I
|
CORETSE_AHBoOiI
)
CORETSE_AHBiloI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBOoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
~
CORETSE_AHBI0oI
&
~
CORETSE_AHBO1oI
)
CORETSE_AHBOoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBiloI
;
end
assign
CORETSE_AHBOlOI
=
CORETSE_AHBO0oI
;
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBI0oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBO1oI
)
CORETSE_AHBI0oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI0oI
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBIoi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIoi
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0oI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBloi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
~
CORETSE_AHBl1oI
)
CORETSE_AHBloi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl1oI
)
CORETSE_AHBloi
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBi0oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1i
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBO1oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO1oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0oI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBI1oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI1oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1i
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBl1oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1oI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBo1oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo1oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiOI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBi1oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi1oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1oI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBOOiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOOiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIII
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBIOiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIOiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOiI
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBiIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOiI
;
end
assign
CORETSE_AHBlOiI
=
CORETSE_AHBIOiI
&
~
CORETSE_AHBiIOI
;
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBO10I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0oI
&
CORETSE_AHBlOo
)
CORETSE_AHBO10I
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBl0oI
&
CORETSE_AHBoOo
)
CORETSE_AHBO10I
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBOOo
or
posedge
CORETSE_AHBilII
)
begin
if
(
CORETSE_AHBilII
)
CORETSE_AHBoOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1oI
)
CORETSE_AHBoOOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
(
CORETSE_AHBl0oI
&
CORETSE_AHBoOo
&
~
CORETSE_AHBi1oI
)
|
(
~
CORETSE_AHBl0oI
&
~
CORETSE_AHBO10I
)
)
CORETSE_AHBoOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
endmodule
