// REVISION    : $Revision: 1.1 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_cnvrxi
(
CORETSE_AHBi010
,
CORETSE_AHBOO1
,
CORETSE_AHBo11
,
CORETSE_AHBO110
,
CORETSE_AHBI110
,
CORETSE_AHBl110
,
CORETSE_AHBo110
,
CORETSE_AHBi110
,
CORETSE_AHBOo10
,
CORETSE_AHBIo10
,
CORETSE_AHBlo10
,
CORETSE_AHBO01
,
CORETSE_AHBol
,
CORETSE_AHBoo10
,
CORETSE_AHBio10
)
;
input
CORETSE_AHBi010
;
input
CORETSE_AHBOO1
;
input
[
1
:
0
]
CORETSE_AHBo11
;
input
[
15
:
0
]
CORETSE_AHBO110
;
input
[
1
:
0
]
CORETSE_AHBI110
;
input
[
1
:
0
]
CORETSE_AHBl110
;
input
CORETSE_AHBo110
;
input
[
3
:
0
]
CORETSE_AHBi110
;
output
[
7
:
0
]
CORETSE_AHBOo10
;
output
CORETSE_AHBIo10
;
output
CORETSE_AHBlo10
;
output
CORETSE_AHBO01
;
output
CORETSE_AHBol
;
output
CORETSE_AHBoo10
;
output
[
3
:
0
]
CORETSE_AHBio10
;
`define CORETSE_AHBIoII  \
# \
1
reg
[
15
:
0
]
CORETSE_AHBOi10
;
reg
[
1
:
0
]
CORETSE_AHBIi10
;
reg
[
1
:
0
]
CORETSE_AHBli10
;
reg
[
1
:
0
]
CORETSE_AHBoi10
;
reg
[
5
:
0
]
CORETSE_AHBii10
;
wire
CORETSE_AHBOOo0
;
reg
[
3
:
0
]
CORETSE_AHBIOo0
;
reg
[
9
:
0
]
CORETSE_AHBlOo0
;
reg
[
9
:
0
]
CORETSE_AHBoOo0
;
reg
[
9
:
0
]
CORETSE_AHBiOo0
;
reg
[
9
:
0
]
CORETSE_AHBOIo0
;
reg
[
9
:
0
]
CORETSE_AHBIIo0
;
reg
[
9
:
0
]
CORETSE_AHBlIo0
;
reg
[
9
:
0
]
CORETSE_AHBoIo0
;
reg
[
9
:
0
]
CORETSE_AHBiIo0
;
reg
[
9
:
0
]
CORETSE_AHBOlo0
;
reg
[
9
:
0
]
CORETSE_AHBIlo0
;
reg
[
9
:
0
]
CORETSE_AHBllo0
;
reg
[
9
:
0
]
CORETSE_AHBolo0
;
reg
[
9
:
0
]
CORETSE_AHBilo0
;
reg
[
9
:
0
]
CORETSE_AHBO0o0
;
reg
[
9
:
0
]
CORETSE_AHBI0o0
;
reg
[
9
:
0
]
CORETSE_AHBl0o0
;
wire
[
9
:
0
]
CORETSE_AHBo0o0
;
wire
CORETSE_AHBi0o0
;
wire
CORETSE_AHBO1o0
;
reg
CORETSE_AHBoo10
;
reg
CORETSE_AHBI1o0
;
reg
[
3
:
0
]
CORETSE_AHBio10
;
wire
CORETSE_AHBl1o0
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOi10
<=
`CORETSE_AHBIoII
16
'h
00
;
else
CORETSE_AHBOi10
<=
`CORETSE_AHBIoII
CORETSE_AHBO110
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIi10
<=
`CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBIi10
<=
`CORETSE_AHBIoII
CORETSE_AHBI110
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoi10
<=
`CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBoi10
<=
`CORETSE_AHBIoII
CORETSE_AHBl110
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBli10
<=
`CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBli10
<=
`CORETSE_AHBIoII
CORETSE_AHBIi10
;
end
assign
CORETSE_AHBl1o0
=
CORETSE_AHBo11
==
2
'b
10
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
6
'h
00
;
else
if
(
CORETSE_AHBl1o0
|
(
(
CORETSE_AHBo11
==
2
'b
01
)
&
(
CORETSE_AHBii10
==
6
'd
4
)
)
|
(
(
CORETSE_AHBo11
==
2
'b
00
)
&
(
CORETSE_AHBii10
==
6
'd
49
)
)
)
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
6
'h
00
;
else
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
CORETSE_AHBii10
+
6
'h
01
;
end
assign
CORETSE_AHBOOo0
=
CORETSE_AHBl1o0
|
(
CORETSE_AHBii10
==
6
'h
02
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIOo0
<=
`CORETSE_AHBIoII
4
'h
0
;
else
if
(
CORETSE_AHBOOo0
)
CORETSE_AHBIOo0
<=
`CORETSE_AHBIoII
CORETSE_AHBIOo0
+
4
'h
1
;
end
assign
CORETSE_AHBO1o0
=
(
(
|
CORETSE_AHBIi10
)
&
CORETSE_AHBOOo0
)
|
(
CORETSE_AHBoo10
&
(
|
CORETSE_AHBIi10
)
)
|
(
~
CORETSE_AHBoo10
&
~
CORETSE_AHBI1o0
&
CORETSE_AHBOOo0
)
;
assign
CORETSE_AHBi0o0
=
(
~
(
|
CORETSE_AHBIi10
)
&
CORETSE_AHBOOo0
)
|
(
CORETSE_AHBoo10
&
CORETSE_AHBI1o0
&
CORETSE_AHBOOo0
)
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoo10
<=
`CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBO1o0
)
CORETSE_AHBoo10
<=
`CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBi0o0
)
CORETSE_AHBoo10
<=
`CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBio10
<=
`CORETSE_AHBIoII
4
'h
0
;
else
if
(
~
CORETSE_AHBoo10
&
CORETSE_AHBO1o0
&
(
CORETSE_AHBo11
==
2
'b
10
)
)
CORETSE_AHBio10
<=
`CORETSE_AHBIoII
CORETSE_AHBIOo0
-
4
'h
1
;
else
if
(
~
CORETSE_AHBoo10
&
CORETSE_AHBO1o0
)
CORETSE_AHBio10
<=
`CORETSE_AHBIoII
CORETSE_AHBIOo0
-
4
'h
6
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBI1o0
<=
`CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBOOo0
)
CORETSE_AHBI1o0
<=
`CORETSE_AHBIoII
CORETSE_AHBoo10
;
end
assign
CORETSE_AHBol
=
|
CORETSE_AHBI110
;
assign
CORETSE_AHBO01
=
|
CORETSE_AHBI110
&
CORETSE_AHBo110
;
assign
CORETSE_AHBo0o0
=
{
10
{
(
CORETSE_AHBi110
==
4
'h
0
)
}
}
&
CORETSE_AHBlOo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
1
)
}
}
&
CORETSE_AHBoOo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
2
)
}
}
&
CORETSE_AHBiOo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
3
)
}
}
&
CORETSE_AHBOIo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
4
)
}
}
&
CORETSE_AHBIIo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
5
)
}
}
&
CORETSE_AHBlIo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
6
)
}
}
&
CORETSE_AHBoIo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
7
)
}
}
&
CORETSE_AHBiIo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
8
)
}
}
&
CORETSE_AHBOlo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
9
)
}
}
&
CORETSE_AHBIlo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
a
)
}
}
&
CORETSE_AHBllo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
b
)
}
}
&
CORETSE_AHBolo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
c
)
}
}
&
CORETSE_AHBilo0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
d
)
}
}
&
CORETSE_AHBO0o0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
e
)
}
}
&
CORETSE_AHBI0o0
|
{
10
{
(
CORETSE_AHBi110
==
4
'h
f
)
}
}
&
CORETSE_AHBl0o0
;
assign
CORETSE_AHBOo10
=
CORETSE_AHBo0o0
[
7
:
0
]
;
assign
CORETSE_AHBIo10
=
CORETSE_AHBo0o0
[
8
]
;
assign
CORETSE_AHBlo10
=
CORETSE_AHBo0o0
[
9
]
;
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlOo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
0
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
0
)
)
)
CORETSE_AHBlOo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoOo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
0
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
1
)
)
)
CORETSE_AHBoOo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiOo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
1
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
2
)
)
)
CORETSE_AHBiOo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOIo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
1
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
3
)
)
)
CORETSE_AHBOIo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIIo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
2
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
4
)
)
)
CORETSE_AHBIIo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBlIo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
2
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
5
)
)
)
CORETSE_AHBlIo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBoIo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
3
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
6
)
)
)
CORETSE_AHBoIo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBiIo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
3
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
7
)
)
)
CORETSE_AHBiIo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBOlo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
4
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
8
)
)
)
CORETSE_AHBOlo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBIlo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
4
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
9
)
)
)
CORETSE_AHBIlo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBllo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
5
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
10
)
)
)
CORETSE_AHBllo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBolo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
5
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
11
)
)
)
CORETSE_AHBolo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBilo0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
6
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
12
)
)
)
CORETSE_AHBilo0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBO0o0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
6
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
13
)
)
)
CORETSE_AHBO0o0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBI0o0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
7
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
14
)
)
)
CORETSE_AHBI0o0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
0
]
,
CORETSE_AHBIi10
[
0
]
,
CORETSE_AHBOi10
[
7
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBOO1
or
posedge
CORETSE_AHBi010
)
begin
if
(
CORETSE_AHBi010
)
CORETSE_AHBl0o0
<=
`CORETSE_AHBIoII
10
'h
000
;
else
if
(
(
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
2
:
0
]
==
3
'd
7
)
)
|
(
~
CORETSE_AHBl1o0
&
(
CORETSE_AHBIOo0
[
3
:
0
]
==
4
'd
15
)
)
)
CORETSE_AHBl0o0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBoi10
[
1
]
,
CORETSE_AHBIi10
[
1
]
,
CORETSE_AHBOi10
[
15
:
8
]
}
;
end
endmodule
