//                        Proprietary and Confidential                          
//                  Copyright (c) 2014 All Rights Reserved                     
// REVISION    : $Revision: 1.7 $                                                  
module
sib_sync_pulse
#
(
parameter
CORETSE_AHBo1IoI
=
0
,
parameter
CORETSE_AHBloloI
=
0
)
(
input
CORETSE_AHBO0I,
input
CORETSE_AHBooloI,
input
CORETSE_AHBioloI,
input
CORETSE_AHBI0I,
input
CORETSE_AHBOiloI,
output
CORETSE_AHBIiloI,
output
CORETSE_AHBliloI
)
;
wire
CORETSE_AHBoiloI
,
CORETSE_AHBiOi1
;
reg
CORETSE_AHBiiloI
,
CORETSE_AHBOO0oI
,
CORETSE_AHBIO0oI
;
wire
CORETSE_AHBlO0oI
,
CORETSE_AHBoO0oI
;
generate
if
(
CORETSE_AHBloloI
==
0
)
begin
:
CORETSE_AHBiO0oI
assign
CORETSE_AHBoiloI
=
CORETSE_AHBiiloI
^
(
!
CORETSE_AHBiOi1
&
CORETSE_AHBioloI
)
;
assign
CORETSE_AHBiOi1
=
CORETSE_AHBlO0oI
^
CORETSE_AHBiiloI
;
assign
CORETSE_AHBliloI
=
CORETSE_AHBlO0oI
^
CORETSE_AHBIO0oI
;
assign
CORETSE_AHBIiloI
=
CORETSE_AHBoO0oI
^
CORETSE_AHBOO0oI
;
sib_sync_2flp
#
(
.CORETSE_AHBlIloI
(
1
)
,
.CORETSE_AHBoIloI
(
CORETSE_AHBo1IoI
)
)
CORETSE_AHBOI0oI
(
.CORETSE_AHBOlloI
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBIlloI
(
CORETSE_AHBO0I
)
,
.CORETSE_AHBllloI
(
CORETSE_AHBOiloI
)
,
.CORETSE_AHBolloI
(
CORETSE_AHBooloI
)
,
.CORETSE_AHBilloI
(
CORETSE_AHBOO0oI
)
,
.CORETSE_AHBO0loI
(
CORETSE_AHBlO0oI
)
)
;
sib_sync_2flp
#
(
.CORETSE_AHBlIloI
(
1
)
,
.CORETSE_AHBoIloI
(
CORETSE_AHBo1IoI
)
)
CORETSE_AHBII0oI
(
.CORETSE_AHBOlloI
(
CORETSE_AHBO0I
)
,
.CORETSE_AHBIlloI
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBllloI
(
CORETSE_AHBooloI
)
,
.CORETSE_AHBolloI
(
CORETSE_AHBOiloI
)
,
.CORETSE_AHBilloI
(
CORETSE_AHBiiloI
)
,
.CORETSE_AHBO0loI
(
CORETSE_AHBoO0oI
)
)
;
always
@
(
posedge
CORETSE_AHBO0I
or
negedge
CORETSE_AHBooloI
)
begin
if
(
!
CORETSE_AHBooloI
)
begin
CORETSE_AHBiiloI
<=
'b
0
;
CORETSE_AHBIO0oI
<=
'b
0
;
end
else
begin
CORETSE_AHBiiloI
<=
CORETSE_AHBoiloI
;
CORETSE_AHBIO0oI
<=
CORETSE_AHBlO0oI
;
end
end
always
@
(
posedge
CORETSE_AHBI0I
or
negedge
CORETSE_AHBOiloI
)
begin
if
(
!
CORETSE_AHBOiloI
)
CORETSE_AHBOO0oI
<=
'b
0
;
else
CORETSE_AHBOO0oI
<=
CORETSE_AHBoO0oI
;
end
end
else
begin
:
CORETSE_AHBlI0oI
assign
CORETSE_AHBIiloI
=
CORETSE_AHBioloI
;
assign
CORETSE_AHBliloI
=
1
'b
1
;
end
endgenerate
endmodule
