// REVISION    : $Revision: 1.20 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
perfn_top
#
(
parameter
CORETSE_AHBoOI
=
0
,
parameter
CORETSE_AHBlOI
=
0
)
(
CORETSE_AHBo111
,
CORETSE_AHBi1Oo
,
CORETSE_AHBiI
,
CORETSE_AHBlI
,
CORETSE_AHBIl
,
CORETSE_AHBol
,
CORETSE_AHBI0Io
,
CORETSE_AHBoo01
,
CORETSE_AHBOOOo
,
CORETSE_AHBio01
,
CORETSE_AHBi0i1
,
CORETSE_AHBO1i1
,
CORETSE_AHBIii1
,
CORETSE_AHBloOo
,
CORETSE_AHBIiIo
,
CORETSE_AHBliIo
,
CORETSE_AHBoiIo
,
CORETSE_AHBlio1
,
CORETSE_AHBIOi1
,
CORETSE_AHBo0o
,
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
,
CORETSE_AHBOIo1
,
CORETSE_AHBiOo1
,
CORETSE_AHBo1o
,
CORETSE_AHBl1o
,
CORETSE_AHBO1o1
,
CORETSE_AHBI1o1
,
CORETSE_AHBl1o1
,
CORETSE_AHBo1o1
,
CORETSE_AHBi1o1
,
CORETSE_AHBlIo1
,
CORETSE_AHBIIo1
,
CORETSE_AHBiI00
,
CORETSE_AHBOl00
)
;
input
CORETSE_AHBo111
,
CORETSE_AHBi1Oo
;
input
CORETSE_AHBiI
;
input
[
7
:
0
]
CORETSE_AHBlI
;
input
CORETSE_AHBIl
;
input
CORETSE_AHBol
;
input
CORETSE_AHBI0Io
;
input
[
1
:
0
]
CORETSE_AHBoo01
;
input
CORETSE_AHBOOOo
,
CORETSE_AHBio01
,
CORETSE_AHBi0i1
;
input
CORETSE_AHBO1i1
;
input
[
7
:
0
]
CORETSE_AHBIii1
;
input
[
15
:
0
]
CORETSE_AHBloOo
;
input
CORETSE_AHBIiIo
,
CORETSE_AHBliIo
,
CORETSE_AHBoiIo
;
input
CORETSE_AHBlio1
;
output
CORETSE_AHBIOi1
;
output
[
7
:
0
]
CORETSE_AHBo0o
;
output
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
;
output
CORETSE_AHBOIo1
,
CORETSE_AHBiOo1
;
output
CORETSE_AHBo1o
;
output
[
32
:
0
]
CORETSE_AHBl1o
;
output
CORETSE_AHBlIo1
;
output
[
8
:
0
]
CORETSE_AHBIIo1
;
output
CORETSE_AHBiI00
,
CORETSE_AHBOl00
;
output
[
7
:
0
]
CORETSE_AHBO1o1
;
output
[
7
:
0
]
CORETSE_AHBI1o1
;
output
CORETSE_AHBl1o1
;
output
CORETSE_AHBo1o1
;
output
CORETSE_AHBi1o1
;
reg
CORETSE_AHBIOi1
;
reg
[
7
:
0
]
CORETSE_AHBo0o
;
reg
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
;
reg
CORETSE_AHBOIo1
,
CORETSE_AHBiOo1
;
reg
CORETSE_AHBo1o
;
reg
[
32
:
0
]
CORETSE_AHBl1o
;
reg
CORETSE_AHBlIo1
;
reg
[
8
:
0
]
CORETSE_AHBIIo1
;
reg
CORETSE_AHBiI00
,
CORETSE_AHBOl00
;
reg
CORETSE_AHBoIlOI
;
wire
CORETSE_AHBiIlOI
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBOllOI
,
CORETSE_AHBIllOI
;
reg
[
7
:
0
]
CORETSE_AHBlllOI
;
reg
CORETSE_AHBollOI
;
reg
CORETSE_AHBillOI
;
wire
[
7
:
0
]
CORETSE_AHBI1IOI
;
reg
[
7
:
0
]
CORETSE_AHBOii0
;
reg
CORETSE_AHBO0lOI
;
wire
CORETSE_AHBI0lOI
;
reg
CORETSE_AHBl0lOI
;
wire
CORETSE_AHBo0lOI
;
reg
CORETSE_AHBi0lOI
,
CORETSE_AHBO1lOI
;
wire
CORETSE_AHBlOi1
;
reg
CORETSE_AHBI1lOI
,
CORETSE_AHBl1lOI
;
wire
CORETSE_AHBo1lOI
;
reg
CORETSE_AHBi1lOI
,
CORETSE_AHBOolOI
;
wire
CORETSE_AHBIolOI
,
CORETSE_AHBlolOI
,
CORETSE_AHBoolOI
,
CORETSE_AHBiolOI
,
CORETSE_AHBOilOI
,
CORETSE_AHBIilOI
;
reg
CORETSE_AHBlilOI
,
CORETSE_AHBoilOI
,
CORETSE_AHBiilOI
,
CORETSE_AHBOO0OI
,
CORETSE_AHBIO0OI
;
wire
CORETSE_AHBlO0OI
;
reg
CORETSE_AHBoO0OI
;
wire
CORETSE_AHBiO0OI
,
CORETSE_AHBOI0OI
;
wire
[
7
:
0
]
CORETSE_AHBII0OI
;
reg
[
7
:
0
]
CORETSE_AHBlI0OI
;
wire
CORETSE_AHBoI0OI
;
wire
CORETSE_AHBiI0OI
,
CORETSE_AHBOl0OI
;
wire
[
15
:
0
]
CORETSE_AHBIl0OI
;
reg
[
15
:
0
]
CORETSE_AHBll0OI
;
wire
CORETSE_AHBol0OI
,
CORETSE_AHBil0OI
,
CORETSE_AHBO00OI
,
CORETSE_AHBI00OI
;
wire
CORETSE_AHBl00OI
,
CORETSE_AHBo00OI
,
CORETSE_AHBi00OI
,
CORETSE_AHBO10OI
;
wire
CORETSE_AHBI10OI
,
CORETSE_AHBl10OI
,
CORETSE_AHBo10OI
;
wire
CORETSE_AHBi10OI
,
CORETSE_AHBOo0OI
;
wire
CORETSE_AHBIo0OI
,
CORETSE_AHBlo0OI
;
wire
[
14
:
0
]
CORETSE_AHBoo0OI
;
reg
[
14
:
0
]
CORETSE_AHBio0OI
;
wire
CORETSE_AHBOi0OI
;
reg
CORETSE_AHBIi0OI
;
wire
CORETSE_AHBli0OI
;
reg
CORETSE_AHBoi0OI
;
wire
CORETSE_AHBii0OI
;
reg
CORETSE_AHBOO1OI
;
wire
CORETSE_AHBIO1OI
,
CORETSE_AHBlO1OI
,
CORETSE_AHBoO1OI
;
reg
CORETSE_AHBiO1OI
,
CORETSE_AHBOI1OI
;
wire
[
7
:
0
]
CORETSE_AHBII1OI
;
reg
[
7
:
0
]
CORETSE_AHBlI1OI
;
wire
CORETSE_AHBoI1OI
,
CORETSE_AHBiI1OI
,
CORETSE_AHBOl1OI
;
reg
CORETSE_AHBIl1OI
,
CORETSE_AHBll1OI
,
CORETSE_AHBol1OI
;
reg
CORETSE_AHBil1OI
;
wire
[
7
:
0
]
CORETSE_AHBO01OI
;
wire
CORETSE_AHBI01OI
,
CORETSE_AHBl01OI
,
CORETSE_AHBo01OI
;
wire
CORETSE_AHBi01OI
,
CORETSE_AHBO11OI
;
wire
CORETSE_AHBI11OI
,
CORETSE_AHBl11OI
,
CORETSE_AHBo11OI
;
reg
CORETSE_AHBil1o
,
CORETSE_AHBol1o
,
CORETSE_AHBO01o
;
wire
[
31
:
0
]
CORETSE_AHBl01o
;
wire
CORETSE_AHBo01o
;
wire
CORETSE_AHBi11OI
;
wire
[
8
:
0
]
CORETSE_AHBOo1OI
;
wire
CORETSE_AHBIo1OI
;
wire
CORETSE_AHBlo1OI
;
wire
CORETSE_AHBoo1OI
,
CORETSE_AHBio1OI
;
wire
[
15
:
0
]
CORETSE_AHBOi1OI
;
reg
[
15
:
0
]
CORETSE_AHBIi1OI
;
wire
CORETSE_AHBli1OI
,
CORETSE_AHBoi1OI
;
wire
CORETSE_AHBii1OI
;
reg
CORETSE_AHBOOoOI
;
wire
CORETSE_AHBIOoOI
;
reg
CORETSE_AHBlOoOI
;
wire
[
15
:
0
]
CORETSE_AHBoOoOI
;
reg
[
15
:
0
]
CORETSE_AHBiOoOI
;
wire
CORETSE_AHBOIoOI
;
reg
CORETSE_AHBIIoOI
;
wire
CORETSE_AHBlIoOI
;
reg
CORETSE_AHBoIoOI
;
wire
CORETSE_AHBiIoOI
;
reg
CORETSE_AHBOloOI
;
wire
CORETSE_AHBIloOI
;
reg
CORETSE_AHBlloOI
;
wire
CORETSE_AHBoloOI
;
reg
CORETSE_AHBiloOI
;
wire
CORETSE_AHBO0oOI
;
reg
CORETSE_AHBI0oOI
;
wire
CORETSE_AHBl0oOI
;
reg
CORETSE_AHBo0oOI
;
reg
CORETSE_AHBi0oOI
;
wire
CORETSE_AHBO1oOI
;
wire
[
32
:
0
]
CORETSE_AHBI1oOI
;
wire
CORETSE_AHBl1oOI
;
assign
CORETSE_AHBO1o1
=
CORETSE_AHBI1IOI
;
assign
CORETSE_AHBI1o1
=
CORETSE_AHBOii0
;
assign
CORETSE_AHBl1o1
=
CORETSE_AHBiolOI
;
assign
CORETSE_AHBo1o1
=
CORETSE_AHBIO0OI
;
assign
CORETSE_AHBi1o1
=
CORETSE_AHBoilOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOllOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOllOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiI
&
~
CORETSE_AHBOI1OI
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIllOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIllOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiI
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBlllOI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlllOI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBlI
[
7
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBollOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBollOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBillOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBillOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOllOI
;
end
assign
CORETSE_AHBI1IOI
[
7
:
0
]
=
{
8
{
~
CORETSE_AHBoo01
[
1
]
}
}
&
{
CORETSE_AHBlllOI
[
3
:
0
]
,
CORETSE_AHBOii0
[
7
:
4
]
}
|
{
8
{
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBlllOI
[
7
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOii0
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOii0
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1IOI
[
7
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBO0lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBO0lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBollOI
;
end
assign
CORETSE_AHBI0lOI
=
~
CORETSE_AHBoo01
[
1
]
&
(
~
CORETSE_AHBlO0OI
|
CORETSE_AHBlO0OI
&
CORETSE_AHBillOI
&
~
CORETSE_AHBl0lOI
)
|
CORETSE_AHBoo01
[
1
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBl0lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBl0lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0lOI
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBi0lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBi0lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0Io
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBO1lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBO1lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0lOI
;
end
assign
CORETSE_AHBlOi1
=
~
CORETSE_AHBio01
&
CORETSE_AHBO1lOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBI1lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBI1lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBl1lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBl1lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1lOI
;
end
assign
CORETSE_AHBo1lOI
=
CORETSE_AHBl1lOI
&
~
CORETSE_AHBio01
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBi1lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBi1lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOOo
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOolOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOolOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1lOI
;
end
assign
CORETSE_AHBl1oOI
=
~
CORETSE_AHBillOI
&
CORETSE_AHBOolOI
|
CORETSE_AHBillOI
&
CORETSE_AHBIOi1
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIOi1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIOi1
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1oOI
;
end
assign
CORETSE_AHBIolOI
=
CORETSE_AHBlilOI
&
CORETSE_AHBillOI
|
CORETSE_AHBoilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
~
CORETSE_AHBoI0OI
|
CORETSE_AHBiilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
~
CORETSE_AHBoI0OI
|
CORETSE_AHBOO0OI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
~
CORETSE_AHBoI0OI
|
CORETSE_AHBIO0OI
&
CORETSE_AHBillOI
&
|
CORETSE_AHBOii0
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBlilOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlilOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIolOI
;
end
assign
CORETSE_AHBlolOI
=
CORETSE_AHBlilOI
&
~
CORETSE_AHBillOI
|
CORETSE_AHBiilOI
&
~
CORETSE_AHBillOI
|
CORETSE_AHBOO0OI
&
~
CORETSE_AHBillOI
|
CORETSE_AHBIO0OI
&
~
CORETSE_AHBillOI
|
CORETSE_AHBoilOI
&
(
~
CORETSE_AHBillOI
|
CORETSE_AHBlOi1
|
~
CORETSE_AHBl0lOI
|
~
CORETSE_AHBIOi1
)
;
assign
CORETSE_AHBIilOI
=
CORETSE_AHBlolOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBoilOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoilOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIilOI
;
end
assign
CORETSE_AHBoolOI
=
CORETSE_AHBoilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
[
6
:
0
]
!=
7
'b
101_0101
&
CORETSE_AHBl0lOI
&
CORETSE_AHBIOi1
|
CORETSE_AHBOO0OI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
[
6
:
0
]
!=
7
'b
101_0101
&
CORETSE_AHBl0lOI
|
CORETSE_AHBiilOI
&
(
CORETSE_AHBillOI
&
CORETSE_AHBOii0
[
6
:
0
]
!=
7
'b
101_0101
&
CORETSE_AHBl0lOI
|
~
CORETSE_AHBl0lOI
)
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBiilOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiilOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoolOI
;
end
assign
CORETSE_AHBiolOI
=
CORETSE_AHBoilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
0101_0101
&
CORETSE_AHBl0lOI
&
CORETSE_AHBIOi1
|
CORETSE_AHBiilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
0101_0101
&
CORETSE_AHBl0lOI
|
CORETSE_AHBOO0OI
&
(
CORETSE_AHBillOI
&
CORETSE_AHBOii0
!=
8
'b
1101_0101
&
CORETSE_AHBl0lOI
|
~
CORETSE_AHBl0lOI
)
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOO0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOO0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiolOI
;
end
assign
CORETSE_AHBlO0OI
=
CORETSE_AHBoilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBIOi1
|
CORETSE_AHBiilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
|
CORETSE_AHBOO0OI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
|
CORETSE_AHBoO0OI
&
~
CORETSE_AHBoilOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBoO0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoO0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO0OI
;
end
assign
CORETSE_AHBOilOI
=
CORETSE_AHBoilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
CORETSE_AHBoI0OI
&
CORETSE_AHBIOi1
|
CORETSE_AHBiilOI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
CORETSE_AHBoI0OI
|
CORETSE_AHBOO0OI
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
CORETSE_AHBoI0OI
|
CORETSE_AHBIO0OI
&
CORETSE_AHBillOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIO0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIO0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOilOI
;
end
assign
CORETSE_AHBiO0OI
=
CORETSE_AHBIO0OI
&
CORETSE_AHBillOI
;
assign
CORETSE_AHBOI0OI
=
~
(
&
CORETSE_AHBlI0OI
[
7
:
0
]
)
&
(
CORETSE_AHBlilOI
|
CORETSE_AHBoilOI
|
CORETSE_AHBiilOI
|
CORETSE_AHBOO0OI
|
CORETSE_AHBIO0OI
&
~
CORETSE_AHBillOI
)
;
assign
CORETSE_AHBII0OI
[
7
:
0
]
=
{
8
{
~
CORETSE_AHBiO0OI
&
CORETSE_AHBOI0OI
}
}
&
CORETSE_AHBlI0OI
[
7
:
0
]
+
1
'b
1
|
{
8
{
~
CORETSE_AHBiO0OI
&
~
CORETSE_AHBOI0OI
}
}
&
CORETSE_AHBlI0OI
[
7
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBlI0OI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlI0OI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBII0OI
[
7
:
0
]
;
end
assign
CORETSE_AHBoI0OI
=
~
CORETSE_AHBoo01
[
1
]
&
(
CORETSE_AHBlI0OI
[
7
:
0
]
>=
(
CORETSE_AHBIii1
[
7
:
2
]
-
1
'b
1
)
)
|
CORETSE_AHBoo01
[
1
]
&
(
CORETSE_AHBlI0OI
[
7
:
0
]
>=
(
CORETSE_AHBIii1
[
7
:
3
]
-
1
'b
1
)
)
;
assign
CORETSE_AHBiI0OI
=
CORETSE_AHBo1o
;
assign
CORETSE_AHBOl0OI
=
~
(
&
CORETSE_AHBll0OI
[
15
:
0
]
)
&
(
CORETSE_AHBIO0OI
&
CORETSE_AHBl0lOI
&
CORETSE_AHBillOI
)
;
assign
CORETSE_AHBIl0OI
[
15
:
0
]
=
{
16
{
~
CORETSE_AHBiI0OI
&
CORETSE_AHBOl0OI
}
}
&
CORETSE_AHBll0OI
[
15
:
0
]
+
1
'b
1
|
{
16
{
~
CORETSE_AHBiI0OI
&
~
CORETSE_AHBOl0OI
}
}
&
CORETSE_AHBll0OI
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBll0OI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBll0OI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl0OI
[
15
:
0
]
;
end
assign
CORETSE_AHBol0OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0000
;
assign
CORETSE_AHBil0OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0001
;
assign
CORETSE_AHBO00OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0002
;
assign
CORETSE_AHBI00OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0003
;
assign
CORETSE_AHBl00OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0004
;
assign
CORETSE_AHBo00OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0005
;
assign
CORETSE_AHBi00OI
=
CORETSE_AHBll0OI
[
15
:
0
]
>
16
'h
0005
;
assign
CORETSE_AHBO10OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0006
;
assign
CORETSE_AHBI10OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
000c
;
assign
CORETSE_AHBl10OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
000d
;
assign
CORETSE_AHBo1oOI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
000e
;
assign
CORETSE_AHBo10OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
000f
;
assign
CORETSE_AHBi10OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0010
;
assign
CORETSE_AHBOo0OI
=
CORETSE_AHBll0OI
[
15
:
0
]
==
16
'h
0011
;
assign
CORETSE_AHBIo0OI
=
~
CORETSE_AHBo1lOI
|
CORETSE_AHBo1o
;
assign
CORETSE_AHBlo0OI
=
CORETSE_AHBo1lOI
;
assign
CORETSE_AHBoo0OI
[
14
:
0
]
=
{
15
{
~
CORETSE_AHBIo0OI
&
CORETSE_AHBlo0OI
}
}
&
CORETSE_AHBio0OI
[
14
:
0
]
+
1
'b
1
|
{
15
{
~
CORETSE_AHBIo0OI
&
~
CORETSE_AHBlo0OI
}
}
&
CORETSE_AHBio0OI
[
14
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBio0OI
[
14
:
0
]
<=
#
CORETSE_AHBIoII
15
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBio0OI
[
14
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0OI
[
14
:
0
]
;
end
assign
CORETSE_AHBOi0OI
=
~
CORETSE_AHBIi0OI
&
CORETSE_AHBo1lOI
&
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBio0OI
[
14
:
0
]
==
15
'h
30D4
|
~
CORETSE_AHBIi0OI
&
CORETSE_AHBo1lOI
&
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBio0OI
[
14
:
0
]
==
15
'h
186A
|
CORETSE_AHBIi0OI
&
~
CORETSE_AHBo1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIi0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIi0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi0OI
;
end
assign
CORETSE_AHBii0OI
=
CORETSE_AHBOI1OI
&
CORETSE_AHBIllOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOO1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOO1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBii0OI
;
end
assign
CORETSE_AHBIO1OI
=
~
CORETSE_AHBiO1OI
&
CORETSE_AHBOO1OI
&
CORETSE_AHBIllOI
|
CORETSE_AHBiO1OI
&
~
CORETSE_AHBo1o
&
~
CORETSE_AHBO1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBiO1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiO1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIO1OI
;
end
assign
CORETSE_AHBoO1OI
=
CORETSE_AHBoo01
[
0
]
&
(
CORETSE_AHBll0OI
[
15
:
0
]
==
CORETSE_AHBloOo
[
15
:
0
]
-
1
)
&
~
CORETSE_AHBO1i1
|
CORETSE_AHBoo01
[
1
]
&
(
CORETSE_AHBll0OI
[
15
:
0
]
==
CORETSE_AHBloOo
[
15
:
0
]
-
3
)
&
~
CORETSE_AHBO1i1
;
assign
CORETSE_AHBlO1OI
=
CORETSE_AHBoO1OI
|
CORETSE_AHBOI1OI
&
CORETSE_AHBIllOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOI1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOI1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO1OI
;
end
assign
CORETSE_AHBII1OI
[
7
:
0
]
=
{
8
{
CORETSE_AHBIO0OI
&
CORETSE_AHBl0lOI
}
}
&
CORETSE_AHBOii0
[
7
:
0
]
|
{
8
{
CORETSE_AHBIO0OI
&
~
CORETSE_AHBl0lOI
}
}
&
CORETSE_AHBo0o
[
7
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBlI1OI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlI1OI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBII1OI
[
7
:
0
]
;
end
assign
CORETSE_AHBoI1OI
=
CORETSE_AHBIO0OI
&
CORETSE_AHBillOI
&
CORETSE_AHBl0lOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIl1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIl1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI1OI
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBil1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBil1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl1OI
;
end
assign
CORETSE_AHBiI1OI
=
CORETSE_AHBIO0OI
&
CORETSE_AHBl0lOI
&
CORETSE_AHBillOI
&
~
CORETSE_AHBIl1OI
&
~
CORETSE_AHBil1OI
&
~
CORETSE_AHBll1OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBll1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBll1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiI1OI
;
end
assign
CORETSE_AHBOl1OI
=
CORETSE_AHBIO0OI
&
CORETSE_AHBl0lOI
&
~
CORETSE_AHBOllOI
&
CORETSE_AHBillOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBol1OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBol1OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOl1OI
;
end
assign
CORETSE_AHBO01OI
[
7
:
0
]
=
{
8
{
~
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBlI1OI
[
7
:
0
]
|
{
8
{
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBII1OI
[
7
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBo0o
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBo0o
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBO01OI
[
7
:
0
]
;
end
assign
CORETSE_AHBI01OI
=
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBIl1OI
|
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBoI1OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBi0o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBi0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBI01OI
;
end
assign
CORETSE_AHBl01OI
=
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBll1OI
|
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBiI1OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBO1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBO1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBl01OI
;
end
assign
CORETSE_AHBo01OI
=
~
CORETSE_AHBoo01
[
1
]
&
(
CORETSE_AHBol1OI
|
CORETSE_AHBIO0OI
&
~
CORETSE_AHBl0lOI
&
~
CORETSE_AHBOllOI
&
CORETSE_AHBillOI
)
|
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOl1OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBI1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBI1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBo01OI
;
end
assign
CORETSE_AHBO11OI
=
CORETSE_AHBii1OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBiOo1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBO11OI
;
end
assign
CORETSE_AHBi01OI
=
1
'b
0
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOIo1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOIo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBi01OI
;
end
assign
CORETSE_AHBI11OI
=
CORETSE_AHBoilOI
&
~
CORETSE_AHBl11OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBil1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBil1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBI11OI
;
end
assign
CORETSE_AHBl11OI
=
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOilOI
&
CORETSE_AHBOllOI
&
~
CORETSE_AHBl0lOI
|
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOilOI
&
CORETSE_AHBOllOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBol1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBol1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBl11OI
;
end
assign
CORETSE_AHBo11OI
=
~
CORETSE_AHBI11OI
&
~
CORETSE_AHBl11OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBO01o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBO01o
<=
#
CORETSE_AHBIoII
CORETSE_AHBo11OI
;
end
pecrc
CORETSE_AHBi1oOI
(
.CORETSE_AHBOl1o
(
CORETSE_AHBo111
)
,
.CORETSE_AHBIl1o
(
CORETSE_AHBlio1
)
,
.CORETSE_AHBll1o
(
CORETSE_AHBOii0
)
,
.CORETSE_AHBol1o
(
CORETSE_AHBol1o
)
,
.CORETSE_AHBil1o
(
CORETSE_AHBil1o
)
,
.CORETSE_AHBO01o
(
CORETSE_AHBO01o
)
,
.CORETSE_AHBI01o
(
CORETSE_AHBi1Oo
)
,
.CORETSE_AHBl01o
(
CORETSE_AHBl01o
)
,
.CORETSE_AHBo01o
(
CORETSE_AHBo01o
)
)
;
assign
CORETSE_AHBi11OI
=
~
CORETSE_AHBlIo1
&
CORETSE_AHBO10OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBlIo1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlIo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBi11OI
;
end
assign
CORETSE_AHBOo1OI
[
8
:
0
]
=
{
9
{
CORETSE_AHBi11OI
}
}
&
CORETSE_AHBl01o
[
31
:
23
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIIo1
[
8
:
0
]
<=
#
CORETSE_AHBIoII
9
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIIo1
[
8
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOo1OI
[
8
:
0
]
;
end
assign
CORETSE_AHBIo1OI
=
CORETSE_AHBol0OI
&
CORETSE_AHBl0lOI
&
CORETSE_AHBOii0
[
0
]
|
~
(
CORETSE_AHBol0OI
&
CORETSE_AHBl0lOI
)
&
CORETSE_AHBOl00
&
!
CORETSE_AHBiI00
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOl00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOl00
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo1OI
;
end
assign
CORETSE_AHBiIlOI
=
CORETSE_AHBol0OI
&
CORETSE_AHBl0lOI
&
(
&
CORETSE_AHBOii0
[
7
:
0
]
)
|
CORETSE_AHBil0OI
&
CORETSE_AHBl0lOI
&
(
&
CORETSE_AHBOii0
[
7
:
0
]
)
&
CORETSE_AHBoIlOI
|
CORETSE_AHBO00OI
&
CORETSE_AHBl0lOI
&
(
&
CORETSE_AHBOii0
[
7
:
0
]
)
&
CORETSE_AHBoIlOI
|
CORETSE_AHBI00OI
&
CORETSE_AHBl0lOI
&
(
&
CORETSE_AHBOii0
[
7
:
0
]
)
&
CORETSE_AHBoIlOI
|
CORETSE_AHBl00OI
&
CORETSE_AHBl0lOI
&
(
&
CORETSE_AHBOii0
[
7
:
0
]
)
&
CORETSE_AHBoIlOI
|
CORETSE_AHBo00OI
&
CORETSE_AHBl0lOI
&
(
&
CORETSE_AHBOii0
[
7
:
0
]
)
&
CORETSE_AHBoIlOI
|
(
CORETSE_AHBi00OI
|
~
CORETSE_AHBl0lOI
)
&
CORETSE_AHBoIlOI
;
assign
CORETSE_AHBlo1OI
=
CORETSE_AHBi00OI
&
CORETSE_AHBoIlOI
|
~
CORETSE_AHBi00OI
&
1
'b
0
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBoIlOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoIlOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIlOI
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBiI00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiI00
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo1OI
;
end
assign
CORETSE_AHBoo1OI
=
CORETSE_AHBI10OI
&
CORETSE_AHBl0lOI
|
CORETSE_AHBi10OI
&
CORETSE_AHBl0lOI
&
CORETSE_AHBOOoOI
;
assign
CORETSE_AHBio1OI
=
CORETSE_AHBl10OI
&
CORETSE_AHBl0lOI
|
CORETSE_AHBOo0OI
&
CORETSE_AHBl0lOI
&
CORETSE_AHBOOoOI
;
assign
CORETSE_AHBOi1OI
[
15
:
0
]
=
{
16
{
CORETSE_AHBoo1OI
}
}
&
{
CORETSE_AHBOii0
[
7
:
0
]
,
CORETSE_AHBIi1OI
[
7
:
0
]
}
|
{
16
{
CORETSE_AHBio1OI
}
}
&
{
CORETSE_AHBIi1OI
[
15
:
8
]
,
CORETSE_AHBOii0
[
7
:
0
]
}
|
{
16
{
~
CORETSE_AHBoo1OI
&
~
CORETSE_AHBio1OI
}
}
&
{
CORETSE_AHBIi1OI
[
15
:
8
]
,
CORETSE_AHBIi1OI
[
7
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIi1OI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIi1OI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi1OI
[
15
:
0
]
;
end
assign
CORETSE_AHBli1OI
=
CORETSE_AHBIi1OI
[
15
:
0
]
>
16
'h
05dc
;
assign
CORETSE_AHBoi1OI
=
(
CORETSE_AHBIi1OI
[
15
:
0
]
>=
16
'h
002e
)
;
assign
CORETSE_AHBii1OI
=
CORETSE_AHBo10OI
&
CORETSE_AHBl0lOI
&
CORETSE_AHBIi1OI
[
15
:
0
]
==
16
'h
8100
|
(
~
CORETSE_AHBo10OI
|
~
CORETSE_AHBl0lOI
)
&
CORETSE_AHBOOoOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOOoOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOOoOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1OI
;
end
assign
CORETSE_AHBli0OI
=
(
CORETSE_AHBll0OI
[
15
:
0
]
>
16
'h
5ee
)
&
(
CORETSE_AHBll0OI
[
15
:
0
]
<
CORETSE_AHBloOo
[
15
:
0
]
)
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBoi0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoi0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBli0OI
;
end
assign
CORETSE_AHBoOoOI
=
{
16
{
~
CORETSE_AHBOOoOI
&
CORETSE_AHBll0OI
>
5
'h
12
}
}
&
(
CORETSE_AHBll0OI
[
15
:
0
]
-
5
'h
11
)
|
{
16
{
CORETSE_AHBOOoOI
&
CORETSE_AHBll0OI
>
5
'h
16
}
}
&
(
CORETSE_AHBll0OI
[
15
:
0
]
-
5
'h
15
)
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBiOoOI
<=
#
CORETSE_AHBIoII
16
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiOoOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOoOI
;
end
assign
CORETSE_AHBOIoOI
=
CORETSE_AHBoi1OI
&
~
CORETSE_AHBli1OI
&
CORETSE_AHBIi1OI
[
15
:
0
]
!=
CORETSE_AHBiOoOI
[
15
:
0
]
&
CORETSE_AHBi0i1
|
~
CORETSE_AHBoi1OI
&
CORETSE_AHBi0i1
&
CORETSE_AHBiOoOI
[
15
:
0
]
>
16
'h
002e
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBIIoOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIIoOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIoOI
;
end
assign
CORETSE_AHBlIoOI
=
~
CORETSE_AHBoIoOI
&
CORETSE_AHBOllOI
&
CORETSE_AHBollOI
|
CORETSE_AHBoIoOI
&
~
CORETSE_AHBo1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBoIoOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoIoOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIoOI
;
end
assign
CORETSE_AHBiIoOI
=
~
CORETSE_AHBOloOI
&
~
CORETSE_AHBOllOI
&
~
CORETSE_AHBO0lOI
&
CORETSE_AHBollOI
&
CORETSE_AHBlllOI
[
7
:
0
]
==
8
'h
0e
|
CORETSE_AHBOloOI
&
~
CORETSE_AHBo1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBOloOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOloOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIoOI
;
end
assign
CORETSE_AHBIloOI
=
~
CORETSE_AHBlloOI
&
~
CORETSE_AHBillOI
&
CORETSE_AHBol0OI
&
CORETSE_AHBoO0OI
&
CORETSE_AHBIO0OI
|
~
CORETSE_AHBlloOI
&
~
CORETSE_AHBillOI
&
CORETSE_AHBol0OI
&
CORETSE_AHBiilOI
&
~
CORETSE_AHBOO0OI
|
~
CORETSE_AHBlloOI
&
~
CORETSE_AHBillOI
&
CORETSE_AHBol0OI
&
CORETSE_AHBOO0OI
&
~
CORETSE_AHBIO0OI
|
CORETSE_AHBlloOI
&
~
CORETSE_AHBo1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBlloOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlloOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIloOI
;
end
assign
CORETSE_AHBoloOI
=
~
CORETSE_AHBiloOI
&
(
CORETSE_AHBoilOI
|
CORETSE_AHBiilOI
|
CORETSE_AHBOO0OI
)
&
CORETSE_AHBillOI
&
CORETSE_AHBOii0
==
8
'b
1101_0101
&
CORETSE_AHBl0lOI
&
~
CORETSE_AHBoI0OI
|
CORETSE_AHBiloOI
&
~
CORETSE_AHBo1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBiloOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiloOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoloOI
;
end
assign
CORETSE_AHBO0oOI
=
~
CORETSE_AHBI0oOI
&
~
CORETSE_AHBOllOI
&
CORETSE_AHBillOI
&
~
CORETSE_AHBl0lOI
&
~
CORETSE_AHBiO1OI
|
CORETSE_AHBI0oOI
&
~
CORETSE_AHBoilOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBI0oOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBI0oOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0oOI
;
end
assign
CORETSE_AHBl0oOI
=
~
CORETSE_AHBo0oOI
&
~
CORETSE_AHBOllOI
&
CORETSE_AHBillOI
&
CORETSE_AHBIO0OI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBo0oOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBo0oOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0oOI
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBi0oOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBi0oOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0oOI
;
end
assign
CORETSE_AHBO1oOI
=
CORETSE_AHBi0oOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBo1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBo1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1oOI
;
end
assign
CORETSE_AHBI1oOI
[
32
]
=
CORETSE_AHBi0oOI
&
CORETSE_AHBiO1OI
|
~
CORETSE_AHBi0oOI
&
CORETSE_AHBl1o
[
32
]
;
assign
CORETSE_AHBI1oOI
[
31
:
28
]
=
{
4
{
CORETSE_AHBi0oOI
}
}
&
{
CORETSE_AHBIi0OI
,
CORETSE_AHBOOoOI
,
CORETSE_AHBoiIo
,
(
CORETSE_AHBliIo
&
~
CORETSE_AHBoIoOI
&
~
CORETSE_AHBo01o
&
(
CORETSE_AHBll0OI
[
15
:
0
]
>=
16
'h
0040
&
CORETSE_AHBll0OI
[
15
:
0
]
<=
16
'h
5dc
)
)
}
|
{
4
{
~
CORETSE_AHBi0oOI
}
}
&
CORETSE_AHBl1o
[
31
:
28
]
;
assign
CORETSE_AHBI1oOI
[
27
:
24
]
=
{
4
{
CORETSE_AHBi0oOI
}
}
&
{
CORETSE_AHBIiIo
,
CORETSE_AHBI0oOI
,
CORETSE_AHBi00OI
&
CORETSE_AHBiI00
,
CORETSE_AHBi00OI
&
CORETSE_AHBOl00
}
|
{
4
{
~
CORETSE_AHBi0oOI
}
}
&
CORETSE_AHBl1o
[
27
:
24
]
;
assign
CORETSE_AHBI1oOI
[
23
:
20
]
=
{
4
{
CORETSE_AHBi0oOI
}
}
&
{
~
CORETSE_AHBoIoOI
&
~
CORETSE_AHBo01o
,
CORETSE_AHBoi0OI
,
CORETSE_AHBIIoOI
,
CORETSE_AHBo01o
}
|
{
4
{
~
CORETSE_AHBi0oOI
}
}
&
CORETSE_AHBl1o
[
23
:
20
]
;
assign
CORETSE_AHBI1oOI
[
19
:
16
]
=
{
4
{
CORETSE_AHBi0oOI
}
}
&
{
CORETSE_AHBoIoOI
,
CORETSE_AHBOloOI
,
CORETSE_AHBlloOI
,
CORETSE_AHBiloOI
}
|
{
4
{
~
CORETSE_AHBi0oOI
}
}
&
CORETSE_AHBl1o
[
19
:
16
]
;
assign
CORETSE_AHBI1oOI
[
15
:
0
]
=
{
16
{
CORETSE_AHBi0oOI
}
}
&
CORETSE_AHBll0OI
[
15
:
0
]
|
{
16
{
~
CORETSE_AHBi0oOI
}
}
&
CORETSE_AHBl1o
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBlio1
)
begin
if
(
CORETSE_AHBlio1
)
CORETSE_AHBl1o
[
32
:
0
]
<=
#
CORETSE_AHBIoII
33
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBl1o
[
32
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1oOI
[
32
:
0
]
;
end
endmodule
