// REVISION    : $Revision: 1.2 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_peanx_top
(
CORETSE_AHBiOO1
,
CORETSE_AHBOo1
,
CORETSE_AHBOIO1
,
CORETSE_AHBIIO1
,
CORETSE_AHBlIO1
,
CORETSE_AHBoIO1
,
CORETSE_AHBiIO1
,
CORETSE_AHBOlO1
,
CORETSE_AHBIlO1
,
CORETSE_AHBllO1
,
CORETSE_AHBolO1
,
CORETSE_AHBilO1
,
CORETSE_AHBO0O1
,
CORETSE_AHBI0O1
,
CORETSE_AHBl0O1
,
CORETSE_AHBo0O1
,
CORETSE_AHBi0O1
,
CORETSE_AHBO1O1
,
CORETSE_AHBI1O1
,
CORETSE_AHBl1O1
,
CORETSE_AHBo1O1
,
CORETSE_AHBi1O1
,
CORETSE_AHBOoO1
,
CORETSE_AHBIoO1
,
CORETSE_AHBloO1
,
CORETSE_AHBooO1
,
CORETSE_AHBioO1
,
CORETSE_AHBOiO1
,
CORETSE_AHBI1i0
)
;
input
CORETSE_AHBiOO1
;
input
CORETSE_AHBOo1
;
input
CORETSE_AHBOIO1
;
input
CORETSE_AHBIIO1
;
input
CORETSE_AHBlIO1
;
input
[
15
:
0
]
CORETSE_AHBoIO1
;
input
CORETSE_AHBiIO1
;
input
CORETSE_AHBOlO1
;
input
[
15
:
0
]
CORETSE_AHBIlO1
;
input
CORETSE_AHBllO1
;
input
[
15
:
0
]
CORETSE_AHBolO1
;
input
CORETSE_AHBilO1
;
input
CORETSE_AHBO0O1
;
input
CORETSE_AHBI0O1
;
input
CORETSE_AHBl0O1
;
input
CORETSE_AHBo0O1
;
input
CORETSE_AHBi0O1
;
input
CORETSE_AHBO1O1
;
input
CORETSE_AHBI1O1
;
output
CORETSE_AHBl1O1
;
output
CORETSE_AHBo1O1
;
output
CORETSE_AHBi1O1
;
output
[
15
:
0
]
CORETSE_AHBOoO1
;
output
[
15
:
0
]
CORETSE_AHBIoO1
;
output
CORETSE_AHBloO1
;
output
CORETSE_AHBooO1
;
output
[
1
:
0
]
CORETSE_AHBioO1
;
output
[
15
:
0
]
CORETSE_AHBOiO1
;
output
[
8
:
0
]
CORETSE_AHBI1i0
;
reg
CORETSE_AHBl1O1
;
reg
CORETSE_AHBo1O1
;
wire
CORETSE_AHBi1O1
;
reg
[
15
:
0
]
CORETSE_AHBOoO1
;
reg
[
15
:
0
]
CORETSE_AHBIoO1
;
reg
CORETSE_AHBloO1
;
reg
CORETSE_AHBooO1
;
reg
[
1
:
0
]
CORETSE_AHBioO1
;
reg
[
15
:
0
]
CORETSE_AHBOiO1
;
parameter
CORETSE_AHBIoII
=
1
;
wire
CORETSE_AHBIiO1
;
wire
CORETSE_AHBliO1
,
CORETSE_AHBoiO1
,
CORETSE_AHBiiO1
,
CORETSE_AHBOOI1
,
CORETSE_AHBIOI1
;
wire
CORETSE_AHBlOI1
,
CORETSE_AHBoOI1
,
CORETSE_AHBiOI1
,
CORETSE_AHBOII1
;
reg
CORETSE_AHBIII1
,
CORETSE_AHBlII1
,
CORETSE_AHBoII1
,
CORETSE_AHBiII1
,
CORETSE_AHBOlI1
;
reg
CORETSE_AHBIlI1
,
CORETSE_AHBllI1
,
CORETSE_AHBolI1
,
CORETSE_AHBilI1
;
wire
CORETSE_AHBO0I1
,
CORETSE_AHBI0I1
;
wire
CORETSE_AHBl0I1
,
CORETSE_AHBo0I1
,
CORETSE_AHBi0I1
;
wire
CORETSE_AHBO1I1
,
CORETSE_AHBI1I1
,
CORETSE_AHBl1I1
,
CORETSE_AHBo1I1
;
wire
CORETSE_AHBi1I1
,
CORETSE_AHBOoI1
,
CORETSE_AHBIoI1
,
CORETSE_AHBloI1
;
reg
CORETSE_AHBooI1
;
reg
[
20
:
0
]
CORETSE_AHBioI1
;
wire
CORETSE_AHBOiI1
,
CORETSE_AHBIiI1
,
CORETSE_AHBliI1
;
reg
CORETSE_AHBoiI1
;
wire
CORETSE_AHBiiI1
;
wire
CORETSE_AHBOOl1
;
wire
CORETSE_AHBIOl1
;
wire
[
15
:
0
]
CORETSE_AHBlOl1
;
wire
[
15
:
0
]
CORETSE_AHBoOl1
;
wire
CORETSE_AHBiOl1
;
reg
CORETSE_AHBOIl1
;
wire
CORETSE_AHBIIl1
;
wire
[
1
:
0
]
CORETSE_AHBlIl1
;
wire
[
15
:
0
]
CORETSE_AHBoIl1
;
wire
CORETSE_AHBiIl1
;
wire
CORETSE_AHBOll1
;
wire
CORETSE_AHBIll1
;
reg
CORETSE_AHBlll1
;
wire
CORETSE_AHBoll1
;
reg
CORETSE_AHBill1
;
wire
CORETSE_AHBO0l1
;
reg
CORETSE_AHBI0l1
;
wire
CORETSE_AHBl0l1
;
reg
CORETSE_AHBo0l1
;
wire
CORETSE_AHBi0l1
;
reg
CORETSE_AHBO1l1
;
wire
[
15
:
0
]
CORETSE_AHBI1l1
;
reg
[
15
:
0
]
CORETSE_AHBl1l1
;
wire
CORETSE_AHBo1l1
;
wire
CORETSE_AHBi1l1
,
CORETSE_AHBOol1
,
CORETSE_AHBIol1
;
wire
[
1
:
0
]
CORETSE_AHBlol1
;
reg
[
1
:
0
]
CORETSE_AHBool1
;
wire
CORETSE_AHBiol1
;
reg
CORETSE_AHBOil1
;
wire
[
15
:
0
]
CORETSE_AHBIil1
;
reg
[
15
:
0
]
CORETSE_AHBlil1
;
wire
CORETSE_AHBoil1
;
wire
CORETSE_AHBiil1
,
CORETSE_AHBOO01
,
CORETSE_AHBIO01
;
wire
[
1
:
0
]
CORETSE_AHBlO01
;
reg
[
1
:
0
]
CORETSE_AHBoO01
;
wire
CORETSE_AHBiO01
;
reg
CORETSE_AHBOI01
;
wire
[
15
:
0
]
CORETSE_AHBII01
;
reg
[
15
:
0
]
CORETSE_AHBlI01
;
wire
CORETSE_AHBoI01
;
reg
CORETSE_AHBiI01
;
wire
[
2
:
0
]
CORETSE_AHBOl01
;
reg
[
2
:
0
]
CORETSE_AHBIl01
;
wire
CORETSE_AHBll01
;
wire
[
20
:
0
]
CORETSE_AHBol01
;
reg
[
20
:
0
]
CORETSE_AHBil01
;
wire
CORETSE_AHBO001
,
CORETSE_AHBI001
;
reg
CORETSE_AHBl001
,
CORETSE_AHBo001
;
wire
CORETSE_AHBi001
;
reg
CORETSE_AHBO101
;
wire
CORETSE_AHBI101
;
reg
CORETSE_AHBl101
;
wire
CORETSE_AHBo101
;
peanx_sync
CORETSE_AHBi101
(
.CORETSE_AHBiOO1
(
CORETSE_AHBiOO1
)
,
.CORETSE_AHBOo1
(
CORETSE_AHBOo1
)
,
.CORETSE_AHBOIO1
(
CORETSE_AHBOIO1
)
,
.CORETSE_AHBIIO1
(
CORETSE_AHBIIO1
)
,
.CORETSE_AHBlIO1
(
CORETSE_AHBlIO1
)
,
.CORETSE_AHBiIO1
(
CORETSE_AHBiIO1
)
,
.CORETSE_AHBOlO1
(
CORETSE_AHBOlO1
)
,
.CORETSE_AHBllO1
(
CORETSE_AHBllO1
)
,
.CORETSE_AHBilO1
(
CORETSE_AHBilO1
)
,
.CORETSE_AHBO0O1
(
CORETSE_AHBO0O1
)
,
.CORETSE_AHBI0O1
(
CORETSE_AHBI0O1
)
,
.CORETSE_AHBl0O1
(
CORETSE_AHBl0O1
)
,
.CORETSE_AHBo0O1
(
CORETSE_AHBo0O1
)
,
.CORETSE_AHBi0O1
(
CORETSE_AHBi0O1
)
,
.CORETSE_AHBO1O1
(
CORETSE_AHBO1O1
)
,
.CORETSE_AHBI1O1
(
CORETSE_AHBI1O1
)
,
.CORETSE_AHBOoI1
(
CORETSE_AHBOoI1
)
,
.CORETSE_AHBIoI1
(
CORETSE_AHBIoI1
)
,
.CORETSE_AHBloI1
(
CORETSE_AHBloI1
)
,
.CORETSE_AHBOiI1
(
CORETSE_AHBOiI1
)
,
.CORETSE_AHBIiI1
(
CORETSE_AHBIiI1
)
,
.CORETSE_AHBO0I1
(
CORETSE_AHBO0I1
)
,
.CORETSE_AHBI0I1
(
CORETSE_AHBI0I1
)
,
.CORETSE_AHBl0I1
(
CORETSE_AHBl0I1
)
,
.CORETSE_AHBo1I1
(
CORETSE_AHBo1I1
)
,
.CORETSE_AHBi1I1
(
CORETSE_AHBi1I1
)
,
.CORETSE_AHBI1I1
(
CORETSE_AHBI1I1
)
,
.CORETSE_AHBl1I1
(
CORETSE_AHBl1I1
)
,
.CORETSE_AHBO1I1
(
CORETSE_AHBO1I1
)
,
.CORETSE_AHBi0I1
(
CORETSE_AHBi0I1
)
,
.CORETSE_AHBo0I1
(
CORETSE_AHBo0I1
)
,
.CORETSE_AHBo101
(
CORETSE_AHBo101
)
)
;
assign
CORETSE_AHBIiO1
=
CORETSE_AHBl0I1
|
CORETSE_AHBooI1
|
CORETSE_AHBlll1
|
(
CORETSE_AHBIIO1
&
(
CORETSE_AHBioO1
!=
2
'b
10
)
)
;
assign
CORETSE_AHBliO1
=
CORETSE_AHBIiO1
|
CORETSE_AHBiII1
&
(
CORETSE_AHBOI01
&
~
CORETSE_AHBoI01
|
CORETSE_AHBOil1
&
CORETSE_AHBoIO1
==
16
'h
0
)
|
CORETSE_AHBOlI1
&
CORETSE_AHBOil1
&
CORETSE_AHBoIO1
==
16
'h
0
|
CORETSE_AHBllI1
&
CORETSE_AHBOil1
&
CORETSE_AHBoIO1
==
16
'h
0
|
CORETSE_AHBolI1
&
CORETSE_AHBOil1
|
CORETSE_AHBIlI1
&
CORETSE_AHBOil1
&
CORETSE_AHBoIO1
==
16
'h
0
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIII1
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBIII1
<=
#
CORETSE_AHBIoII
CORETSE_AHBliO1
;
end
assign
CORETSE_AHBoiO1
=
CORETSE_AHBIII1
&
~
CORETSE_AHBIiO1
&
CORETSE_AHBO0I1
|
CORETSE_AHBlII1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBo001
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBlII1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlII1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiO1
;
end
assign
CORETSE_AHBOII1
=
CORETSE_AHBIII1
&
~
CORETSE_AHBIiO1
&
~
CORETSE_AHBO0I1
|
CORETSE_AHBilI1
&
~
CORETSE_AHBIiO1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBilI1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBilI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOII1
;
end
assign
CORETSE_AHBiiO1
=
CORETSE_AHBlII1
&
~
CORETSE_AHBIiO1
&
CORETSE_AHBo001
|
CORETSE_AHBoII1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBOil1
&
CORETSE_AHBoIO1
!=
16
'h
0
&
CORETSE_AHBoiI1
|
CORETSE_AHBIoI1
&
CORETSE_AHBi0I1
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBoII1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoII1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiO1
;
end
assign
CORETSE_AHBOOI1
=
CORETSE_AHBoII1
&
CORETSE_AHBOil1
&
|
CORETSE_AHBoIO1
|
CORETSE_AHBIlI1
&
CORETSE_AHBOil1
&
|
CORETSE_AHBoIO1
&
(
CORETSE_AHBO1l1
^
CORETSE_AHBoIO1
[
11
]
)
&
CORETSE_AHBoiI1
|
CORETSE_AHBiII1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBOI01
|
CORETSE_AHBOil1
&
~|
CORETSE_AHBoIO1
&
CORETSE_AHBoiI1
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBiII1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiII1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOI1
;
end
assign
CORETSE_AHBIOI1
=
CORETSE_AHBiII1
&
CORETSE_AHBOI01
&
CORETSE_AHBoI01
|
CORETSE_AHBOlI1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBOil1
&
~|
CORETSE_AHBoIO1
|
CORETSE_AHBoOI1
|
CORETSE_AHBlOI1
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOlI1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOlI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOI1
;
end
assign
CORETSE_AHBoOI1
=
CORETSE_AHBOlI1
&
CORETSE_AHBo001
&
(
(
~
CORETSE_AHBIlO1
[
15
]
&
~
CORETSE_AHBo1I1
|
~
CORETSE_AHBOoO1
[
15
]
)
|
CORETSE_AHBIlO1
[
15
]
&
~
CORETSE_AHBo1I1
&
CORETSE_AHBOoO1
[
15
]
&
~
CORETSE_AHBOiO1
[
15
]
&
~
CORETSE_AHBill1
)
&
(
~
CORETSE_AHBOil1
|
(
|
CORETSE_AHBoIO1
)
)
|
CORETSE_AHBllI1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBOil1
&
~|
CORETSE_AHBoIO1
|
CORETSE_AHBo001
&
CORETSE_AHBll01
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBllI1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBllI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOI1
;
end
assign
CORETSE_AHBiOI1
=
~
CORETSE_AHBolI1
&
CORETSE_AHBllI1
&
CORETSE_AHBo001
&
CORETSE_AHBll01
|
~
CORETSE_AHBolI1
&
CORETSE_AHBoII1
&
CORETSE_AHBIoI1
&
CORETSE_AHBi0I1
|
CORETSE_AHBolI1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBOil1
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBolI1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBolI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOI1
;
end
assign
CORETSE_AHBI1i0
=
{
CORETSE_AHBolI1
,
CORETSE_AHBllI1
,
CORETSE_AHBOlI1
,
CORETSE_AHBIlI1
,
CORETSE_AHBiII1
,
CORETSE_AHBoII1
,
CORETSE_AHBlII1
,
CORETSE_AHBIII1
,
CORETSE_AHBilI1
}
;
assign
CORETSE_AHBlOI1
=
CORETSE_AHBOlI1
&
CORETSE_AHBo001
&
CORETSE_AHBIlO1
[
15
]
&
~
CORETSE_AHBo1I1
&
CORETSE_AHBOoO1
[
15
]
&
CORETSE_AHBl1I1
&
(
CORETSE_AHBOiO1
[
15
]
|
CORETSE_AHBill1
)
&
(
~
CORETSE_AHBOil1
|
(
|
CORETSE_AHBoIO1
)
)
|
CORETSE_AHBIlI1
&
~
(
CORETSE_AHBIiO1
|
CORETSE_AHBOil1
&
~|
CORETSE_AHBoIO1
|
CORETSE_AHBOil1
&
(
CORETSE_AHBO1l1
^
CORETSE_AHBoIO1
[
11
]
)
&
|
CORETSE_AHBoIO1
&
CORETSE_AHBoiI1
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIlI1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIlI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOI1
;
end
assign
CORETSE_AHBliI1
=
CORETSE_AHBOiI1
&
~
CORETSE_AHBIiI1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBoiI1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoiI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBliI1
;
end
assign
CORETSE_AHBIll1
=
CORETSE_AHBO0I1
&
~
CORETSE_AHBI0I1
|
~
CORETSE_AHBO0I1
&
CORETSE_AHBI0I1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBlll1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlll1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIll1
;
end
assign
CORETSE_AHBiiI1
=
~
CORETSE_AHBloO1
&
CORETSE_AHBOlI1
|
CORETSE_AHBloO1
&
~
(
CORETSE_AHBIII1
|
CORETSE_AHBI1I1
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBloO1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBloO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiI1
;
end
assign
CORETSE_AHBoll1
=
CORETSE_AHBl101
&
CORETSE_AHBoIO1
[
15
]
|
~
CORETSE_AHBl101
&
CORETSE_AHBill1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBill1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBill1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoll1
;
end
assign
CORETSE_AHBOOl1
=
~
CORETSE_AHBl1O1
&
CORETSE_AHBolI1
|
CORETSE_AHBl1O1
&
~
CORETSE_AHBIII1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl1O1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1O1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOl1
;
end
assign
CORETSE_AHBIIl1
=
|
CORETSE_AHBoIO1
[
13
:
12
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo1O1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo1O1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIl1
;
end
assign
CORETSE_AHBlIl1
[
1
:
0
]
=
{
2
{
CORETSE_AHBIII1
&
CORETSE_AHBO0I1
|
CORETSE_AHBlII1
}
}
&
2
'b
00
|
{
2
{
CORETSE_AHBIII1
&
~
CORETSE_AHBO0I1
|
CORETSE_AHBllI1
}
}
&
2
'b
01
|
{
2
{
CORETSE_AHBilI1
|
CORETSE_AHBolI1
}
}
&
2
'b
10
|
{
2
{
~
(
CORETSE_AHBIII1
|
CORETSE_AHBlII1
|
CORETSE_AHBllI1
|
CORETSE_AHBilI1
|
CORETSE_AHBolI1
)
}
}
&
CORETSE_AHBioO1
[
1
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBioO1
[
1
:
0
]
<=
#
CORETSE_AHBIoII
2
'b
00
;
else
CORETSE_AHBioO1
[
1
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIl1
[
1
:
0
]
;
end
assign
CORETSE_AHBi001
=
CORETSE_AHBlOI1
&
~
CORETSE_AHBIlI1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBO101
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBO101
<=
#
CORETSE_AHBIoII
CORETSE_AHBi001
;
end
assign
CORETSE_AHBiIl1
=
(
CORETSE_AHBIII1
&
CORETSE_AHBO0I1
)
|
CORETSE_AHBlII1
;
assign
CORETSE_AHBOll1
=
~
(
CORETSE_AHBiIl1
|
CORETSE_AHBoII1
&
~
CORETSE_AHBOil1
&
~
CORETSE_AHBo1I1
|
CORETSE_AHBoII1
&
CORETSE_AHBOil1
&
CORETSE_AHBOI01
&
|
CORETSE_AHBoIO1
|
CORETSE_AHBiII1
|
CORETSE_AHBO101
&
~
CORETSE_AHBi1I1
|
CORETSE_AHBO1I1
)
;
assign
CORETSE_AHBoIl1
=
{
16
{
CORETSE_AHBoII1
&
~
CORETSE_AHBOil1
&
~
CORETSE_AHBo1I1
&
~
CORETSE_AHBiIl1
}
}
&
{
CORETSE_AHBIlO1
[
15
]
,
1
'b
0
,
CORETSE_AHBIlO1
[
13
:
0
]
}
|
{
16
{
(
CORETSE_AHBoII1
&
CORETSE_AHBOil1
&
CORETSE_AHBOI01
&
|
CORETSE_AHBoIO1
&
~
CORETSE_AHBiIl1
)
|
(
CORETSE_AHBiII1
&
~
CORETSE_AHBiIl1
)
}
}
&
{
CORETSE_AHBOiO1
[
15
]
,
1
'b
1
,
CORETSE_AHBOiO1
[
13
:
0
]
}
|
{
16
{
CORETSE_AHBO101
&
~
CORETSE_AHBi1I1
&
~
CORETSE_AHBiIl1
}
}
&
{
CORETSE_AHBolO1
[
15
]
,
1
'b
0
,
CORETSE_AHBolO1
[
13
:
12
]
,
CORETSE_AHBo0l1
,
CORETSE_AHBolO1
[
10
:
0
]
}
|
{
16
{
CORETSE_AHBO1I1
&
~
CORETSE_AHBiIl1
}
}
&
CORETSE_AHBIlO1
|
{
16
{
CORETSE_AHBOll1
}
}
&
CORETSE_AHBOiO1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOiO1
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBOiO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIl1
;
end
assign
CORETSE_AHBIOl1
=
CORETSE_AHBlII1
|
CORETSE_AHBIlI1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBooO1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBooO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOl1
;
end
assign
CORETSE_AHBi1O1
=
CORETSE_AHBolI1
|
CORETSE_AHBilI1
;
wire
CORETSE_AHBOo01
;
assign
CORETSE_AHBOo01
=
CORETSE_AHBIOI1
&
~
CORETSE_AHBOlI1
;
assign
CORETSE_AHBi0l1
=
(
(
CORETSE_AHBOo01
&
CORETSE_AHBoIO1
[
11
]
)
|
(
~
CORETSE_AHBOo01
&
CORETSE_AHBO1l1
)
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBO1l1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO1l1
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0l1
;
end
assign
CORETSE_AHBl0l1
=
CORETSE_AHBoII1
&
CORETSE_AHBIlO1
[
11
]
&
~
CORETSE_AHBo1I1
|
CORETSE_AHBI0l1
&
~
CORETSE_AHBo0l1
|
~
CORETSE_AHBI0l1
&
~
(
CORETSE_AHBoII1
&
~
CORETSE_AHBo1I1
)
&
CORETSE_AHBo0l1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo0l1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo0l1
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0l1
;
end
assign
CORETSE_AHBO0l1
=
CORETSE_AHBIOI1
&
~
CORETSE_AHBOlI1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBI0l1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI0l1
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0l1
;
end
assign
CORETSE_AHBI1l1
=
{
16
{
CORETSE_AHBliI1
&
CORETSE_AHBool1
==
2
'h
0
}
}
&
CORETSE_AHBoIO1
[
15
:
0
]
|
{
16
{
~
CORETSE_AHBliI1
|
CORETSE_AHBool1
!=
2
'h
0
}
}
&
CORETSE_AHBl1l1
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl1l1
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBl1l1
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1l1
;
end
assign
CORETSE_AHBo1l1
=
(
{
CORETSE_AHBl1l1
[
15
]
,
CORETSE_AHBl1l1
[
13
:
0
]
}
==
{
CORETSE_AHBoIO1
[
15
]
,
CORETSE_AHBoIO1
[
13
:
0
]
}
)
&
CORETSE_AHBoIO1
!=
16
'h
0
;
assign
CORETSE_AHBi1l1
=
CORETSE_AHBIoI1
|
CORETSE_AHBloI1
|
CORETSE_AHBliI1
&
(
|
CORETSE_AHBool1
)
&
~
CORETSE_AHBo1l1
|
CORETSE_AHBIII1
|
CORETSE_AHBlII1
;
assign
CORETSE_AHBOol1
=
CORETSE_AHBliI1
&
(
~|
CORETSE_AHBool1
)
;
assign
CORETSE_AHBIol1
=
CORETSE_AHBliI1
&
(
^
CORETSE_AHBool1
)
&
CORETSE_AHBo1l1
;
assign
CORETSE_AHBlol1
[
1
:
0
]
=
{
2
{
CORETSE_AHBi1l1
}
}
&
2
'h
0
|
{
2
{
CORETSE_AHBOol1
}
}
&
2
'h
1
|
{
2
{
CORETSE_AHBIol1
}
}
&
CORETSE_AHBool1
[
1
:
0
]
+
2
'h
1
|
{
2
{
~
CORETSE_AHBi1l1
&
~
CORETSE_AHBOol1
&
~
CORETSE_AHBIol1
}
}
&
CORETSE_AHBool1
[
1
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBool1
<=
#
CORETSE_AHBIoII
2
'h
0
;
else
CORETSE_AHBool1
<=
#
CORETSE_AHBIoII
CORETSE_AHBlol1
;
end
assign
CORETSE_AHBiol1
=
CORETSE_AHBlol1
==
2
'h
3
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOil1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOil1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiol1
;
end
assign
CORETSE_AHBIil1
=
{
16
{
CORETSE_AHBliI1
&
CORETSE_AHBoO01
==
2
'h
0
}
}
&
CORETSE_AHBoIO1
[
15
:
0
]
|
{
16
{
~
CORETSE_AHBliI1
|
CORETSE_AHBoO01
!=
2
'h
0
}
}
&
CORETSE_AHBlil1
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBlil1
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBlil1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIil1
;
end
assign
CORETSE_AHBoil1
=
CORETSE_AHBlil1
[
15
:
0
]
==
CORETSE_AHBoIO1
[
15
:
0
]
;
assign
CORETSE_AHBiil1
=
CORETSE_AHBIoI1
|
CORETSE_AHBloI1
|
~
CORETSE_AHBoIO1
[
14
]
|
CORETSE_AHBliI1
&
CORETSE_AHBoO01
>
2
'h
0
&
CORETSE_AHBoIO1
[
14
]
&
~
CORETSE_AHBoil1
|
CORETSE_AHBlII1
;
assign
CORETSE_AHBOO01
=
~
CORETSE_AHBiil1
&
CORETSE_AHBliI1
&
~|
CORETSE_AHBoO01
&
CORETSE_AHBoIO1
[
14
]
;
assign
CORETSE_AHBIO01
=
CORETSE_AHBliI1
&
(
^
CORETSE_AHBoO01
)
&
CORETSE_AHBlil1
[
14
]
&
CORETSE_AHBoIO1
[
14
]
&
CORETSE_AHBoil1
;
assign
CORETSE_AHBlO01
=
{
2
{
CORETSE_AHBiil1
}
}
&
2
'h
0
|
{
2
{
CORETSE_AHBOO01
}
}
&
2
'h
1
|
{
2
{
CORETSE_AHBIO01
}
}
&
CORETSE_AHBoO01
+
2
'h
1
|
{
2
{
~
CORETSE_AHBiil1
&
~
CORETSE_AHBOO01
&
~
CORETSE_AHBIO01
}
}
&
CORETSE_AHBoO01
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBoO01
[
1
:
0
]
<=
#
CORETSE_AHBIoII
2
'h
0
;
else
CORETSE_AHBoO01
[
1
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO01
[
1
:
0
]
;
end
assign
CORETSE_AHBiO01
=
CORETSE_AHBlO01
==
2
'h
3
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOI01
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOI01
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO01
;
end
assign
CORETSE_AHBII01
=
{
16
{
CORETSE_AHBoII1
&
CORETSE_AHBool1
==
2
'h
3
|
CORETSE_AHBIlI1
&
CORETSE_AHBool1
==
2
'h
3
}
}
&
CORETSE_AHBl1l1
|
{
16
{
~
(
CORETSE_AHBoII1
&
CORETSE_AHBool1
==
2
'h
3
|
CORETSE_AHBIlI1
&
CORETSE_AHBool1
==
2
'h
3
)
}
}
&
CORETSE_AHBlI01
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBlI01
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBlI01
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBII01
[
15
:
0
]
;
end
assign
CORETSE_AHBoI01
=
CORETSE_AHBOI01
&
{
CORETSE_AHBl1l1
[
15
]
,
CORETSE_AHBl1l1
[
13
:
0
]
}
==
{
CORETSE_AHBlI01
[
15
]
,
CORETSE_AHBlI01
[
13
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBiI01
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBiI01
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI01
;
end
assign
CORETSE_AHBOl01
=
{
3
{
CORETSE_AHBliI1
|
CORETSE_AHBloI1
}
}
&
3
'h
0
|
{
3
{
CORETSE_AHBIoI1
&
~&
CORETSE_AHBIl01
}
}
&
CORETSE_AHBIl01
[
2
:
0
]
+
3
'h
1
|
{
3
{
CORETSE_AHBIoI1
&
(
&
CORETSE_AHBIl01
)
}
}
&
CORETSE_AHBIl01
[
2
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIl01
[
2
:
0
]
<=
#
CORETSE_AHBIoII
3
'h
0
;
else
CORETSE_AHBIl01
[
2
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOl01
[
2
:
0
]
;
end
assign
CORETSE_AHBll01
=
CORETSE_AHBIl01
[
2
:
1
]
==
2
'h
3
;
assign
CORETSE_AHBO001
=
CORETSE_AHBoiO1
&
~
CORETSE_AHBlII1
|
CORETSE_AHBIOI1
&
~
CORETSE_AHBOlI1
|
CORETSE_AHBoOI1
&
~
CORETSE_AHBllI1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl001
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBl001
<=
#
CORETSE_AHBIoII
CORETSE_AHBO001
;
end
assign
CORETSE_AHBI001
=
CORETSE_AHBil01
[
20
:
0
]
==
21
'h
1
|
CORETSE_AHBo001
&
~
CORETSE_AHBO001
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo001
<=
#
CORETSE_AHBIoII
1
'h
1
;
else
CORETSE_AHBo001
<=
#
CORETSE_AHBIoII
CORETSE_AHBI001
;
end
assign
CORETSE_AHBol01
[
20
:
0
]
=
{
21
{
CORETSE_AHBl001
&
~
CORETSE_AHBo0I1
&
~
CORETSE_AHBo101
}
}
&
21
'd
200000
|
{
21
{
CORETSE_AHBl001
&
~
CORETSE_AHBo0I1
&
CORETSE_AHBo101
}
}
&
21
'h
13_12D0
|
{
21
{
CORETSE_AHBl001
&
CORETSE_AHBo0I1
}
}
&
21
'h
00_0040
|
{
21
{
~
CORETSE_AHBl001
&
|
CORETSE_AHBil01
[
20
:
0
]
}
}
&
CORETSE_AHBil01
-
21
'h
1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBil01
[
20
:
0
]
<=
#
CORETSE_AHBIoII
21
'h
0
;
else
CORETSE_AHBil01
[
20
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBol01
[
20
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBioI1
[
20
:
0
]
<=
#
CORETSE_AHBIoII
21
'h
0
;
else
if
(
CORETSE_AHBOoI1
&
~
CORETSE_AHBo0I1
)
CORETSE_AHBioI1
[
20
:
0
]
<=
#
CORETSE_AHBIoII
21
'h
13_12D0
;
else
if
(
CORETSE_AHBOoI1
&
CORETSE_AHBo0I1
)
CORETSE_AHBioI1
[
20
:
0
]
<=
#
CORETSE_AHBIoII
21
'h
00_0040
;
else
if
(
|
CORETSE_AHBioI1
[
20
:
0
]
)
CORETSE_AHBioI1
[
20
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBioI1
-
21
'h
1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBooI1
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBooI1
<=
#
CORETSE_AHBIoII
(
~
CORETSE_AHBOoI1
&
~
(
|
CORETSE_AHBioI1
[
20
:
0
]
)
)
;
end
assign
CORETSE_AHBI101
=
CORETSE_AHBIOI1
&
~
CORETSE_AHBOlI1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl101
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBl101
<=
#
CORETSE_AHBIoII
CORETSE_AHBI101
;
end
assign
CORETSE_AHBiOl1
=
~
CORETSE_AHBOIl1
&
CORETSE_AHBIlI1
|
CORETSE_AHBOIl1
&
~
CORETSE_AHBIII1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOIl1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOIl1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOl1
;
end
assign
CORETSE_AHBlOl1
=
{
16
{
~
CORETSE_AHBOIl1
&
CORETSE_AHBl101
}
}
&
CORETSE_AHBoIO1
[
15
:
0
]
|
{
16
{
~
(
~
CORETSE_AHBOIl1
&
CORETSE_AHBl101
)
}
}
&
CORETSE_AHBOoO1
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOoO1
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBOoO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOl1
[
15
:
0
]
;
end
assign
CORETSE_AHBoOl1
=
{
16
{
CORETSE_AHBOIl1
&
CORETSE_AHBl101
}
}
&
CORETSE_AHBoIO1
[
15
:
0
]
|
{
16
{
~
(
CORETSE_AHBOIl1
&
CORETSE_AHBl101
)
}
}
&
CORETSE_AHBIoO1
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIoO1
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBIoO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOl1
[
15
:
0
]
;
end
endmodule
