// VERSION     : $Revision: 1.1 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
pecrc
(
CORETSE_AHBOl1o
,
CORETSE_AHBIl1o
,
CORETSE_AHBll1o
,
CORETSE_AHBol1o
,
CORETSE_AHBil1o
,
CORETSE_AHBO01o
,
CORETSE_AHBI01o
,
CORETSE_AHBl01o
,
CORETSE_AHBo01o
)
;
input
CORETSE_AHBOl1o
,
CORETSE_AHBIl1o
;
input
[
7
:
0
]
CORETSE_AHBll1o
;
input
CORETSE_AHBol1o
;
input
CORETSE_AHBil1o
,
CORETSE_AHBO01o
;
input
CORETSE_AHBI01o
;
output
[
31
:
0
]
CORETSE_AHBl01o
;
output
CORETSE_AHBo01o
;
reg
[
31
:
0
]
CORETSE_AHBl01o
;
wire
CORETSE_AHBo01o
;
parameter
CORETSE_AHBIoII
=
1
;
wire
[
7
:
0
]
CORETSE_AHBi01o
;
wire
[
31
:
0
]
CORETSE_AHBO11o
;
reg
[
31
:
0
]
CORETSE_AHBI11o
;
assign
CORETSE_AHBi01o
[
0
]
=
CORETSE_AHBl01o
[
31
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
0
]
)
;
assign
CORETSE_AHBi01o
[
1
]
=
CORETSE_AHBl01o
[
30
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
1
]
)
;
assign
CORETSE_AHBi01o
[
2
]
=
CORETSE_AHBl01o
[
29
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
2
]
)
;
assign
CORETSE_AHBi01o
[
3
]
=
CORETSE_AHBl01o
[
28
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
3
]
)
;
assign
CORETSE_AHBi01o
[
4
]
=
CORETSE_AHBl01o
[
27
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
4
]
)
;
assign
CORETSE_AHBi01o
[
5
]
=
CORETSE_AHBl01o
[
26
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
5
]
)
;
assign
CORETSE_AHBi01o
[
6
]
=
CORETSE_AHBl01o
[
25
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
6
]
)
;
assign
CORETSE_AHBi01o
[
7
]
=
CORETSE_AHBl01o
[
24
]
^
(
CORETSE_AHBol1o
&
CORETSE_AHBll1o
[
7
]
)
;
assign
CORETSE_AHBO11o
[
31
]
=
CORETSE_AHBl01o
[
23
]
^
CORETSE_AHBi01o
[
2
]
;
assign
CORETSE_AHBO11o
[
30
]
=
CORETSE_AHBl01o
[
22
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
3
]
;
assign
CORETSE_AHBO11o
[
29
]
=
CORETSE_AHBl01o
[
21
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
4
]
;
assign
CORETSE_AHBO11o
[
28
]
=
CORETSE_AHBl01o
[
20
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
5
]
;
assign
CORETSE_AHBO11o
[
27
]
=
CORETSE_AHBl01o
[
19
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
26
]
=
CORETSE_AHBl01o
[
18
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
25
]
=
CORETSE_AHBl01o
[
17
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
;
assign
CORETSE_AHBO11o
[
24
]
=
CORETSE_AHBl01o
[
16
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
23
]
=
CORETSE_AHBl01o
[
15
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
22
]
=
CORETSE_AHBl01o
[
14
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
21
]
=
CORETSE_AHBl01o
[
13
]
^
CORETSE_AHBi01o
[
2
]
;
assign
CORETSE_AHBO11o
[
20
]
=
CORETSE_AHBl01o
[
12
]
^
CORETSE_AHBi01o
[
3
]
;
assign
CORETSE_AHBO11o
[
19
]
=
CORETSE_AHBl01o
[
11
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
4
]
;
assign
CORETSE_AHBO11o
[
18
]
=
CORETSE_AHBl01o
[
10
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
5
]
;
assign
CORETSE_AHBO11o
[
17
]
=
CORETSE_AHBl01o
[
9
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
16
]
=
CORETSE_AHBl01o
[
8
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
15
]
=
CORETSE_AHBl01o
[
7
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
;
assign
CORETSE_AHBO11o
[
14
]
=
CORETSE_AHBl01o
[
6
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
;
assign
CORETSE_AHBO11o
[
13
]
=
CORETSE_AHBl01o
[
5
]
^
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
12
]
=
CORETSE_AHBl01o
[
4
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
11
]
=
CORETSE_AHBl01o
[
3
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
10
]
=
CORETSE_AHBl01o
[
2
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
9
]
=
CORETSE_AHBl01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
8
]
=
CORETSE_AHBl01o
[
0
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
7
]
=
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
6
]
=
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
5
]
=
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
2
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
4
]
=
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
3
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
3
]
=
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
4
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
;
assign
CORETSE_AHBO11o
[
2
]
=
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
5
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
1
]
=
CORETSE_AHBi01o
[
0
]
^
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
6
]
^
CORETSE_AHBi01o
[
7
]
;
assign
CORETSE_AHBO11o
[
0
]
=
CORETSE_AHBi01o
[
1
]
^
CORETSE_AHBi01o
[
7
]
;
always
@
(
CORETSE_AHBil1o
or
CORETSE_AHBol1o
or
CORETSE_AHBO01o
or
CORETSE_AHBO11o
or
CORETSE_AHBl01o
)
begin
case
(
1
'b
1
)
CORETSE_AHBil1o
:
CORETSE_AHBI11o
=
32
'h
ffff_ffff
;
CORETSE_AHBol1o
:
CORETSE_AHBI11o
=
CORETSE_AHBO11o
[
31
:
0
]
;
CORETSE_AHBO01o
:
CORETSE_AHBI11o
=
CORETSE_AHBl01o
[
31
:
0
]
;
default
:
CORETSE_AHBI11o
=
32
'h
0000_0000
;
endcase
end
always
@
(
posedge
CORETSE_AHBOl1o
or
posedge
CORETSE_AHBIl1o
)
begin
if
(
CORETSE_AHBIl1o
)
CORETSE_AHBl01o
[
31
:
0
]
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
if
(
CORETSE_AHBI01o
)
CORETSE_AHBl01o
[
31
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBI11o
[
31
:
0
]
;
end
assign
CORETSE_AHBo01o
=
CORETSE_AHBl01o
[
31
:
0
]
!=
32
'b
11000111000001001101110101111011
;
endmodule
