//                     Proprietary and Confidential
// REVISION    : $Revision: $
`include "include.v"
module
ptp_tfp
(
input
CORETSE_AHBOI01I,
input
CORETSE_AHBII01I,
input
CORETSE_AHBlOo0I,
input
CORETSE_AHBlI01I,
input
CORETSE_AHBoI01I,
input
[
1
:
0
]
CORETSE_AHBoIo0I,
input
[
7
:
0
]
CORETSE_AHBiI01I,
input
[
7
:
0
]
CORETSE_AHBOl01I,
input
CORETSE_AHBi1O1I,
input
CORETSE_AHBIl01I,
input
CORETSE_AHBoOo0I,
input
[
79
:
0
]
CORETSE_AHBll01I,
input
CORETSE_AHBol01I,
input
CORETSE_AHBil01I,
output
CORETSE_AHBO001I,
output
[
15
:
0
]
CORETSE_AHBIlo0I,
output
[
79
:
0
]
CORETSE_AHBllo0I,
output
[
3
:
0
]
CORETSE_AHBolo0I,
output
CORETSE_AHBI001I,
output
CORETSE_AHBl001I,
output
[
15
:
0
]
CORETSE_AHBo001I,
output
CORETSE_AHBi001I,
output
CORETSE_AHBO101I,
output
CORETSE_AHBI101I
)
;
reg
[
15
:
0
]
CORETSE_AHBO0o0I
;
wire
[
15
:
0
]
CORETSE_AHBI0o0I
;
reg
[
15
:
0
]
CORETSE_AHBl0o0I
;
wire
[
15
:
0
]
CORETSE_AHBo0o0I
;
wire
[
5
:
0
]
CORETSE_AHBi0o0I
;
wire
CORETSE_AHBIo1II
;
wire
CORETSE_AHBl101I
;
reg
[
3
:
0
]
CORETSE_AHBO1o0I
;
wire
[
3
:
0
]
CORETSE_AHBI1o0I
;
reg
[
7
:
0
]
msg_qu [11 : 0]
;
wire
[
7
:
0
]
msg_qu_c [11 : 0]
;
reg
CORETSE_AHBo101I
;
wire
CORETSE_AHBi101I
;
wire
CORETSE_AHBOo01I
;
reg
CORETSE_AHBIo01I
;
reg
CORETSE_AHBlo01I
;
wire
CORETSE_AHBoo01I
;
wire
CORETSE_AHBio01I
;
wire
CORETSE_AHBOi01I
;
wire
CORETSE_AHBIi01I
;
wire
CORETSE_AHBli01I
;
reg
CORETSE_AHBi1o0I
;
wire
CORETSE_AHBOoo0I
;
reg
CORETSE_AHBoi01I
;
wire
CORETSE_AHBii01I
;
wire
CORETSE_AHBOO11I
;
reg
[
15
:
0
]
CORETSE_AHBIO11I
;
wire
[
15
:
0
]
CORETSE_AHBlO11I
;
reg
CORETSE_AHBooo0I
;
reg
CORETSE_AHBioo0I
;
wire
[
16
:
0
]
CORETSE_AHBoO11I
;
wire
[
16
:
0
]
CORETSE_AHBiO11I
;
wire
[
17
:
0
]
CORETSE_AHBOI11I
;
wire
[
18
:
0
]
CORETSE_AHBII11I
;
reg
[
18
:
0
]
CORETSE_AHBlI11I
;
wire
[
18
:
0
]
CORETSE_AHBoI11I
;
wire
[
19
:
0
]
CORETSE_AHBiI11I
;
wire
CORETSE_AHBOl11I
;
wire
CORETSE_AHBIl11I
;
wire
CORETSE_AHBll11I
;
wire
CORETSE_AHBol11I
;
reg
CORETSE_AHBil11I
;
reg
CORETSE_AHBO011I
;
reg
CORETSE_AHBI011I
;
reg
CORETSE_AHBl011I
;
reg
CORETSE_AHBo011I
;
reg
CORETSE_AHBi011I
;
reg
CORETSE_AHBO111I
;
wire
CORETSE_AHBI111I
;
reg
CORETSE_AHBl111I
;
wire
CORETSE_AHBo111I
;
reg
CORETSE_AHBi111I
;
wire
CORETSE_AHBOo11I
;
reg
CORETSE_AHBIo11I
;
wire
CORETSE_AHBlo11I
;
reg
CORETSE_AHBoo11I
;
wire
CORETSE_AHBio11I
;
reg
CORETSE_AHBOi11I
;
wire
CORETSE_AHBIi11I
;
reg
CORETSE_AHBli11I
;
wire
CORETSE_AHBoi11I
;
reg
CORETSE_AHBii11I
;
wire
CORETSE_AHBOOo1I
;
reg
CORETSE_AHBIOo1I
;
wire
CORETSE_AHBlOo1I
;
reg
CORETSE_AHBoOo1I
;
wire
CORETSE_AHBiOo1I
;
reg
CORETSE_AHBOIo1I
;
wire
CORETSE_AHBIIo1I
;
reg
CORETSE_AHBlIo1I
;
wire
CORETSE_AHBoIo1I
;
reg
CORETSE_AHBiIo1I
;
wire
CORETSE_AHBOlo1I
;
reg
CORETSE_AHBIlo1I
;
wire
CORETSE_AHBllo1I
;
reg
CORETSE_AHBolo1I
;
wire
CORETSE_AHBilo1I
;
wire
CORETSE_AHBooi0I
;
wire
CORETSE_AHBioi0I
;
wire
CORETSE_AHBOii0I
;
wire
CORETSE_AHBO0o1I
;
reg
CORETSE_AHBI0o1I
;
reg
CORETSE_AHBl0o1I
;
wire
CORETSE_AHBOIO1I
;
reg
CORETSE_AHBIIO1I
;
reg
CORETSE_AHBOo1II
;
wire
CORETSE_AHBoIO1I
;
reg
CORETSE_AHBlIO1I
;
reg
CORETSE_AHBo0o1I
;
reg
CORETSE_AHBo1llI
;
wire
CORETSE_AHBi0o1I
;
reg
CORETSE_AHBO1o1I
;
reg
CORETSE_AHBI1o1I
;
wire
CORETSE_AHBl1o1I
;
reg
CORETSE_AHBilI1I
;
reg
CORETSE_AHBo1o1I
;
wire
[
1
:
0
]
CORETSE_AHBoo01
;
reg
[
7
:
0
]
CORETSE_AHBi1o1I
;
reg
[
7
:
0
]
CORETSE_AHBOoo1I
;
wire
CORETSE_AHBIoo1I
;
reg
CORETSE_AHBloo1I
;
wire
[
7
:
0
]
CORETSE_AHBIl0lI
;
wire
[
7
:
0
]
CORETSE_AHBiOIlI
;
assign
CORETSE_AHBO001I
=
CORETSE_AHBlo01I
;
assign
CORETSE_AHBolo0I
=
CORETSE_AHBO1o0I
;
assign
CORETSE_AHBI001I
=
CORETSE_AHBo101I
;
assign
CORETSE_AHBl001I
=
CORETSE_AHBl101I
;
assign
CORETSE_AHBi001I
=
CORETSE_AHBO111I
;
assign
CORETSE_AHBo001I
=
(
~
(
CORETSE_AHBiI11I
[
19
:
16
]
+
CORETSE_AHBiI11I
[
15
:
0
]
)
)
;
assign
CORETSE_AHBI101I
=
(
CORETSE_AHBIO11I
==
16
'b
0
)
;
assign
CORETSE_AHBllo0I
=
{
msg_qu
[
11
]
,
msg_qu
[
10
]
,
msg_qu
[
9
]
,
msg_qu
[
8
]
,
msg_qu
[
7
]
,
msg_qu
[
6
]
,
msg_qu
[
5
]
,
msg_qu
[
4
]
,
msg_qu
[
3
]
,
msg_qu
[
2
]
}
;
assign
CORETSE_AHBIlo0I
=
{
msg_qu
[
1
]
,
msg_qu
[
0
]
}
;
assign
CORETSE_AHBO101I
=
CORETSE_AHBIIO1I
;
assign
CORETSE_AHBIl0lI
=
CORETSE_AHBi1o1I
;
assign
CORETSE_AHBiOIlI
=
CORETSE_AHBOoo1I
;
assign
CORETSE_AHBoo01
=
CORETSE_AHBoIo0I
;
assign
CORETSE_AHBO0o1I
=
CORETSE_AHBII01I
|
CORETSE_AHBlOo0I
;
assign
CORETSE_AHBi0o0I
=
{
CORETSE_AHBiOIlI
[
3
:
0
]
,
2
'b
00
}
-
2
'b
10
;
assign
CORETSE_AHBi101I
=
~
CORETSE_AHBI011I
&
(
~
CORETSE_AHBo1llI
&
CORETSE_AHBOo01I
|
~
CORETSE_AHBo1llI
&
~
CORETSE_AHBOo01I
&
CORETSE_AHBo101I
)
;
assign
CORETSE_AHBl101I
=
~
CORETSE_AHBo1llI
&
CORETSE_AHBIo1II
;
assign
CORETSE_AHBii01I
=
~
CORETSE_AHBo1llI
&
CORETSE_AHBOO11I
;
assign
CORETSE_AHBI111I
=
~
CORETSE_AHBo011I
&
(
CORETSE_AHBoi01I
|
(
~
CORETSE_AHBoi01I
&
CORETSE_AHBi011I
)
)
;
assign
CORETSE_AHBi0o1I
=
CORETSE_AHBo0o1I
|
CORETSE_AHBoI01I
;
assign
CORETSE_AHBl1o1I
=
CORETSE_AHBi1O1I
|
CORETSE_AHBilI1I
;
assign
CORETSE_AHBIoo1I
=
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBilI1I
|
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBo1o1I
;
assign
CORETSE_AHBOIO1I
=
CORETSE_AHBoo01
[
1
]
|
~
CORETSE_AHBoo01
[
1
]
&
(
CORETSE_AHBlIO1I
&
~
CORETSE_AHBOo1II
)
;
assign
CORETSE_AHBoIO1I
=
~
CORETSE_AHBI1o1I
&
(
CORETSE_AHBi1O1I
|
(
~
CORETSE_AHBi1O1I
&
CORETSE_AHBlIO1I
)
)
;
assign
CORETSE_AHBo111I
=
CORETSE_AHBo1llI
|
(
CORETSE_AHBl111I
&
~
(
CORETSE_AHBioo0I
&
CORETSE_AHBloo1I
)
|
CORETSE_AHBii11I
&
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
8
&&
CORETSE_AHBiOIlI
!=
8
'h
11
)
|
CORETSE_AHBIOo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
&&
CORETSE_AHBiOIlI
!=
8
'h
11
)
|
CORETSE_AHBIlo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
2
&&
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
!=
16
'h
013F
)
|
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
0
)
&
(
(
CORETSE_AHBiOIlI
[
3
]
|
CORETSE_AHBiOIlI
[
2
]
)
==
1
'b
1
)
|
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
6
&&
(
~
CORETSE_AHBiOIlI
[
1
]
!=
CORETSE_AHBIl01I
)
)
|
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1F
&&
!
CORETSE_AHBil11I
)
|
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
2B
)
|
(
!
CORETSE_AHBOo11I
&
!
CORETSE_AHBlo11I
&
!
CORETSE_AHBio11I
&
!
CORETSE_AHBIi11I
&
!
CORETSE_AHBoi11I
&
!
CORETSE_AHBOOo1I
&
!
CORETSE_AHBlOo1I
&
!
CORETSE_AHBiOo1I
&
!
CORETSE_AHBIIo1I
&
!
CORETSE_AHBoIo1I
&
!
CORETSE_AHBOlo1I
&
!
CORETSE_AHBllo1I
&
!
CORETSE_AHBilo1I
)
)
;
assign
CORETSE_AHBOo11I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBl111I
&
CORETSE_AHBioo0I
&
CORETSE_AHBloo1I
|
CORETSE_AHBi111I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
A
)
)
;
assign
CORETSE_AHBlo11I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBi111I
&
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
A
)
)
;
assign
CORETSE_AHBio11I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIo11I
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
8100
)
|
CORETSE_AHBOi11I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
8100
)
|
CORETSE_AHBoo11I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
;
assign
CORETSE_AHBIi11I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIo11I
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
88A8
)
|
CORETSE_AHBOi11I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
88A8
)
|
CORETSE_AHBOi11I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
;
assign
CORETSE_AHBoi11I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIo11I
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
8847
||
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
8848
)
|
CORETSE_AHBoo11I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
8847
||
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
8848
)
|
CORETSE_AHBli11I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
;
assign
CORETSE_AHBOOo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBli11I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
&
(
CORETSE_AHBiOIlI
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBiOIlI
[
3
:
0
]
>
4
'h
4
)
|
CORETSE_AHBoOo1I
&
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
&
(
CORETSE_AHBiOIlI
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBiOIlI
[
3
:
0
]
>
4
'h
4
)
|
CORETSE_AHBii11I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
8
&&
CORETSE_AHBiOIlI
!=
8
'h
11
)
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
;
assign
CORETSE_AHBlOo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBli11I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
&
(
CORETSE_AHBiOIlI
[
7
:
4
]
==
4
'h
6
)
|
CORETSE_AHBOIo1I
&
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
|
CORETSE_AHBIOo1I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
;
assign
CORETSE_AHBiOo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIo11I
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
0800
)
|
CORETSE_AHBoo11I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
0800
)
|
CORETSE_AHBoOo1I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
;
assign
CORETSE_AHBIIo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIo11I
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
86DD
)
|
CORETSE_AHBoo11I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
86DD
)
|
CORETSE_AHBOIo1I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
;
assign
CORETSE_AHBoIo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIo11I
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
88F7
)
|
CORETSE_AHBoo11I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
==
16
'h
88F7
)
)
;
assign
CORETSE_AHBOlo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBIOo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
&&
CORETSE_AHBiOIlI
==
8
'h
11
)
|
CORETSE_AHBiIo1I
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
;
assign
CORETSE_AHBllo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBii11I
&
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
|
CORETSE_AHBiIo1I
&
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
|
CORETSE_AHBIlo1I
&
~
(
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
2
&&
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
!=
16
'h
013F
)
)
&
~
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
)
;
assign
CORETSE_AHBilo1I
=
!
CORETSE_AHBo1llI
&
(
CORETSE_AHBlIo1I
|
CORETSE_AHBIlo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
|
CORETSE_AHBolo1I
&
!
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
6
&&
(
~
CORETSE_AHBiOIlI
[
1
]
!=
CORETSE_AHBIl01I
)
)
&
!
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1F
&&
!
CORETSE_AHBil11I
)
&
!
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
2B
)
&
!
(
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
0
)
&
(
(
CORETSE_AHBiOIlI
[
2
]
|
CORETSE_AHBiOIlI
[
3
]
)
==
1
'b
1
)
)
)
;
assign
CORETSE_AHBI1o0I
=
{
4
{
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
0
)
}
}
&
CORETSE_AHBiOIlI
[
3
:
0
]
|
{
4
{
~
(
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
0
)
)
}
}
&
CORETSE_AHBO1o0I
;
assign
CORETSE_AHBIl11I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1
)
&
(
CORETSE_AHBO1o0I
==
4
'h
0
)
&
CORETSE_AHBIl01I
;
assign
CORETSE_AHBIo1II
=
CORETSE_AHBIlo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
&
(
CORETSE_AHBIl0lI
[
3
:
0
]
==
4
'h
0
)
&
CORETSE_AHBIl01I
;
assign
CORETSE_AHBOl11I
=
CORETSE_AHBIlo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
6
)
;
assign
CORETSE_AHBOo01I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
6
&&
(
~
CORETSE_AHBiOIlI
[
1
]
!=
CORETSE_AHBIl01I
)
)
;
assign
CORETSE_AHBOO11I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1F
)
;
assign
CORETSE_AHBll11I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
6
&&
(
~
CORETSE_AHBiOIlI
[
1
]
!=
CORETSE_AHBIl01I
)
)
|
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1F
&&
!
CORETSE_AHBil11I
)
|
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
2B
)
;
assign
CORETSE_AHBOi01I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
2b
)
;
assign
CORETSE_AHBio01I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
21
)
;
assign
CORETSE_AHBIi01I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
13
)
;
assign
CORETSE_AHBli01I
=
CORETSE_AHBolo1I
&
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1F
)
;
assign
CORETSE_AHBI0o0I
=
{
16
{
~
CORETSE_AHBo1llI
}
}
&
(
{
16
{
(
CORETSE_AHBi111I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
A
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBOi11I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBoo11I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBli11I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBoOo1I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBOIo1I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBiIo1I
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBii11I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
8
&&
CORETSE_AHBiOIlI
!=
8
'h
11
)
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBIOo1I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBIlo1I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
2
&&
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
!=
16
'h
013F
)
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBolo1I
&
!
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
6
&&
(
~
CORETSE_AHBiOIlI
[
1
]
!=
CORETSE_AHBIl01I
)
)
&
!
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
1F
&&
!
CORETSE_AHBil11I
)
&
!
(
CORETSE_AHBO0o0I
[
5
:
0
]
==
6
'h
2B
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
)
;
assign
CORETSE_AHBooi0I
=
CORETSE_AHBli11I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
&
(
CORETSE_AHBiOIlI
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBiOIlI
[
3
:
0
]
>
4
'h
4
)
;
assign
CORETSE_AHBioi0I
=
CORETSE_AHBoOo1I
&
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
&
(
CORETSE_AHBiOIlI
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBiOIlI
[
3
:
0
]
>
4
'h
4
)
;
assign
CORETSE_AHBOii0I
=
CORETSE_AHBIOo1I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
3
)
;
assign
CORETSE_AHBo0o0I
=
{
16
{
CORETSE_AHBooi0I
}
}
&
{
10
'b
0
,
CORETSE_AHBi0o0I
}
|
{
16
{
CORETSE_AHBioi0I
}
}
&
{
10
'b
0
,
CORETSE_AHBi0o0I
}
|
{
16
{
CORETSE_AHBOii0I
}
}
&
(
16
'h
28
-
16
'h
8
)
|
{
16
{
~
(
CORETSE_AHBooi0I
|
CORETSE_AHBioi0I
|
CORETSE_AHBOii0I
)
}
}
&
CORETSE_AHBl0o0I
;
assign
CORETSE_AHBoo01I
=
~
CORETSE_AHBOi01I
&
~
CORETSE_AHBo1llI
&
(
CORETSE_AHBio01I
|
~
CORETSE_AHBio01I
&
CORETSE_AHBIo01I
)
;
assign
CORETSE_AHBOoo0I
=
~
CORETSE_AHBli01I
&
~
CORETSE_AHBo1llI
&
(
CORETSE_AHBIi01I
|
(
~
CORETSE_AHBIi01I
&
CORETSE_AHBi1o0I
)
)
;
assign
CORETSE_AHBol11I
=
~
CORETSE_AHBll11I
&
~
CORETSE_AHBo1llI
&
(
CORETSE_AHBIl11I
|
(
~
CORETSE_AHBIl11I
&
CORETSE_AHBil11I
)
)
;
assign
msg_qu_c
[
0
]
=
(
{
8
{
CORETSE_AHBi1o0I
}
}
&
CORETSE_AHBiOIlI
)
|
(
{
8
{
~
CORETSE_AHBi1o0I
}
}
&
msg_qu
[
0
]
)
;
generate
genvar
CORETSE_AHBOloI
;
for
(
CORETSE_AHBOloI
=
1
;
CORETSE_AHBOloI
<
12
;
CORETSE_AHBOloI
=
CORETSE_AHBOloI
+
1
)
begin
:
CORETSE_AHBooo1I
assign
msg_qu_c
[
CORETSE_AHBOloI
]
=
(
{
8
{
CORETSE_AHBi1o0I
}
}
&
msg_qu
[
CORETSE_AHBOloI
-
1
]
)
|
(
{
8
{
~
CORETSE_AHBi1o0I
}
}
&
msg_qu
[
CORETSE_AHBOloI
]
)
;
end
endgenerate
assign
CORETSE_AHBlO11I
=
{
16
{
CORETSE_AHBOl11I
}
}
&
(
~
{
CORETSE_AHBiOIlI
,
CORETSE_AHBIl0lI
}
)
|
{
16
{
~
CORETSE_AHBOl11I
}
}
&
CORETSE_AHBIO11I
;
assign
CORETSE_AHBoO11I
=
CORETSE_AHBll01I
[
15
:
0
]
+
CORETSE_AHBll01I
[
31
:
16
]
;
assign
CORETSE_AHBiO11I
=
CORETSE_AHBll01I
[
47
:
32
]
+
CORETSE_AHBll01I
[
63
:
48
]
;
assign
CORETSE_AHBOI11I
=
CORETSE_AHBoO11I
+
CORETSE_AHBiO11I
;
assign
CORETSE_AHBII11I
=
CORETSE_AHBOI11I
+
CORETSE_AHBll01I
[
79
:
64
]
;
assign
CORETSE_AHBoI11I
=
{
19
{
CORETSE_AHBOl11I
}
}
&
CORETSE_AHBII11I
|
{
19
{
~
CORETSE_AHBOl11I
}
}
&
CORETSE_AHBII11I
;
assign
CORETSE_AHBiI11I
=
CORETSE_AHBlI11I
+
CORETSE_AHBIO11I
;
always
@
(
posedge
CORETSE_AHBOI01I
or
posedge
CORETSE_AHBl0o1I
)
begin
if
(
CORETSE_AHBl0o1I
)
begin
CORETSE_AHBooo0I
<=
1
'b
0
;
CORETSE_AHBioo0I
<=
1
'b
0
;
CORETSE_AHBO011I
<=
1
'b
0
;
CORETSE_AHBI011I
<=
1
'b
0
;
CORETSE_AHBl011I
<=
1
'b
0
;
CORETSE_AHBo011I
<=
1
'b
0
;
CORETSE_AHBi011I
<=
1
'b
0
;
CORETSE_AHBO111I
<=
1
'b
0
;
CORETSE_AHBo0o1I
<=
1
'b
0
;
CORETSE_AHBo1llI
<=
1
'b
0
;
CORETSE_AHBO1o1I
<=
1
'b
0
;
CORETSE_AHBI1o1I
<=
1
'b
0
;
CORETSE_AHBlIO1I
<=
1
'b
0
;
CORETSE_AHBIIO1I
<=
1
'b
0
;
CORETSE_AHBO0o0I
<=
16
'b
0
;
CORETSE_AHBl0o0I
<=
16
'b
0
;
CORETSE_AHBO1o0I
<=
4
'b
0
;
CORETSE_AHBo101I
<=
1
'b
0
;
CORETSE_AHBi1o0I
<=
1
'b
0
;
msg_qu
[
0
]
<=
8
'b
0
;
msg_qu
[
1
]
<=
8
'b
0
;
msg_qu
[
2
]
<=
8
'b
0
;
msg_qu
[
3
]
<=
8
'b
0
;
msg_qu
[
4
]
<=
8
'b
0
;
msg_qu
[
5
]
<=
8
'b
0
;
msg_qu
[
6
]
<=
8
'b
0
;
msg_qu
[
7
]
<=
8
'b
0
;
msg_qu
[
8
]
<=
8
'b
0
;
msg_qu
[
9
]
<=
8
'b
0
;
msg_qu
[
10
]
<=
8
'b
0
;
msg_qu
[
11
]
<=
8
'b
0
;
CORETSE_AHBIo01I
<=
1
'b
0
;
CORETSE_AHBlo01I
<=
1
'b
0
;
CORETSE_AHBoi01I
<=
1
'b
0
;
CORETSE_AHBlI11I
<=
19
'b
0
;
CORETSE_AHBil11I
<=
1
'b
0
;
CORETSE_AHBIO11I
<=
16
'b
1
;
CORETSE_AHBl111I
<=
1
'b
1
;
CORETSE_AHBi111I
<=
1
'b
0
;
CORETSE_AHBIo11I
<=
1
'b
0
;
CORETSE_AHBoo11I
<=
1
'b
0
;
CORETSE_AHBOi11I
<=
1
'b
0
;
CORETSE_AHBli11I
<=
1
'b
0
;
CORETSE_AHBii11I
<=
1
'b
0
;
CORETSE_AHBIOo1I
<=
1
'b
0
;
CORETSE_AHBoOo1I
<=
1
'b
0
;
CORETSE_AHBOIo1I
<=
1
'b
0
;
CORETSE_AHBlIo1I
<=
1
'b
0
;
CORETSE_AHBiIo1I
<=
1
'b
0
;
CORETSE_AHBIlo1I
<=
1
'b
0
;
CORETSE_AHBolo1I
<=
1
'b
0
;
CORETSE_AHBilI1I
<=
1
'b
0
;
CORETSE_AHBo1o1I
<=
1
'b
0
;
CORETSE_AHBi1o1I
<=
8
'b
0
;
CORETSE_AHBOoo1I
<=
8
'b
0
;
CORETSE_AHBloo1I
<=
1
'b
0
;
CORETSE_AHBOo1II
<=
1
'b
0
;
end
else
begin
CORETSE_AHBooo0I
<=
CORETSE_AHBoOo0I
;
CORETSE_AHBioo0I
<=
CORETSE_AHBooo0I
;
CORETSE_AHBO011I
<=
CORETSE_AHBol01I
;
CORETSE_AHBI011I
<=
CORETSE_AHBO011I
;
CORETSE_AHBl011I
<=
CORETSE_AHBil01I
;
CORETSE_AHBo011I
<=
CORETSE_AHBl011I
;
CORETSE_AHBi011I
<=
CORETSE_AHBI111I
;
CORETSE_AHBO111I
<=
CORETSE_AHBi011I
;
CORETSE_AHBo0o1I
<=
CORETSE_AHBoI01I
;
CORETSE_AHBo1llI
<=
CORETSE_AHBi0o1I
;
CORETSE_AHBO1o1I
<=
CORETSE_AHBo1llI
;
CORETSE_AHBI1o1I
<=
CORETSE_AHBO1o1I
;
CORETSE_AHBlIO1I
<=
CORETSE_AHBoIO1I
;
CORETSE_AHBOo1II
<=
CORETSE_AHBOIO1I
;
CORETSE_AHBIIO1I
<=
CORETSE_AHBOo1II
;
CORETSE_AHBi1o1I
<=
CORETSE_AHBOl01I
;
CORETSE_AHBOoo1I
<=
CORETSE_AHBiI01I
;
CORETSE_AHBloo1I
<=
CORETSE_AHBIoo1I
;
CORETSE_AHBilI1I
<=
CORETSE_AHBi1O1I
;
CORETSE_AHBo1o1I
<=
CORETSE_AHBl1o1I
;
CORETSE_AHBlo01I
<=
CORETSE_AHBIo01I
;
if
(
CORETSE_AHBlI01I
&&
CORETSE_AHBIIO1I
)
begin
CORETSE_AHBO0o0I
<=
CORETSE_AHBI0o0I
;
CORETSE_AHBl0o0I
<=
CORETSE_AHBo0o0I
;
CORETSE_AHBO1o0I
<=
CORETSE_AHBI1o0I
;
CORETSE_AHBo101I
<=
CORETSE_AHBi101I
;
CORETSE_AHBi1o0I
<=
CORETSE_AHBOoo0I
;
msg_qu
[
0
]
<=
msg_qu_c
[
0
]
;
msg_qu
[
1
]
<=
msg_qu_c
[
1
]
;
msg_qu
[
2
]
<=
msg_qu_c
[
2
]
;
msg_qu
[
3
]
<=
msg_qu_c
[
3
]
;
msg_qu
[
4
]
<=
msg_qu_c
[
4
]
;
msg_qu
[
5
]
<=
msg_qu_c
[
5
]
;
msg_qu
[
6
]
<=
msg_qu_c
[
6
]
;
msg_qu
[
7
]
<=
msg_qu_c
[
7
]
;
msg_qu
[
8
]
<=
msg_qu_c
[
8
]
;
msg_qu
[
9
]
<=
msg_qu_c
[
9
]
;
msg_qu
[
10
]
<=
msg_qu_c
[
10
]
;
msg_qu
[
11
]
<=
msg_qu_c
[
11
]
;
CORETSE_AHBIo01I
<=
CORETSE_AHBoo01I
;
CORETSE_AHBoi01I
<=
CORETSE_AHBii01I
;
CORETSE_AHBlI11I
<=
CORETSE_AHBoI11I
;
CORETSE_AHBil11I
<=
CORETSE_AHBol11I
;
CORETSE_AHBIO11I
<=
CORETSE_AHBlO11I
;
CORETSE_AHBl111I
<=
CORETSE_AHBo111I
;
CORETSE_AHBi111I
<=
CORETSE_AHBOo11I
;
CORETSE_AHBIo11I
<=
CORETSE_AHBlo11I
;
CORETSE_AHBoo11I
<=
CORETSE_AHBio11I
;
CORETSE_AHBOi11I
<=
CORETSE_AHBIi11I
;
CORETSE_AHBli11I
<=
CORETSE_AHBoi11I
;
CORETSE_AHBii11I
<=
CORETSE_AHBOOo1I
;
CORETSE_AHBIOo1I
<=
CORETSE_AHBlOo1I
;
CORETSE_AHBoOo1I
<=
CORETSE_AHBiOo1I
;
CORETSE_AHBOIo1I
<=
CORETSE_AHBIIo1I
;
CORETSE_AHBlIo1I
<=
CORETSE_AHBoIo1I
;
CORETSE_AHBiIo1I
<=
CORETSE_AHBOlo1I
;
CORETSE_AHBIlo1I
<=
CORETSE_AHBllo1I
;
CORETSE_AHBolo1I
<=
CORETSE_AHBilo1I
;
end
end
end
always
@
(
posedge
CORETSE_AHBOI01I
or
posedge
CORETSE_AHBO0o1I
)
begin
if
(
CORETSE_AHBO0o1I
)
begin
CORETSE_AHBI0o1I
<=
1
'b
1
;
CORETSE_AHBl0o1I
<=
1
'b
1
;
end
else
begin
CORETSE_AHBI0o1I
<=
1
'b
0
;
CORETSE_AHBl0o1I
<=
CORETSE_AHBI0o1I
;
end
end
endmodule
