//               centralization improves synthesis and layout development 
// REVISION    : $Revision: 1.2 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxfif_clkrst
(
CORETSE_AHBIi0
,
CORETSE_AHBoo1
,
CORETSE_AHBoi0
,
CORETSE_AHBii0
,
CORETSE_AHBOOo
,
CORETSE_AHBOlo
,
CORETSE_AHBioOI
,
CORETSE_AHBOiOI
,
CORETSE_AHBIiOI
,
CORETSE_AHBliOI
,
CORETSE_AHBoiOI
,
CORETSE_AHBilII
,
CORETSE_AHBO0II
,
CORETSE_AHBI0II
,
CORETSE_AHBl0II
,
CORETSE_AHBo0II
)
;
input
CORETSE_AHBIi0
;
input
CORETSE_AHBoo1
;
input
CORETSE_AHBoi0
;
input
CORETSE_AHBii0
;
input
CORETSE_AHBOOo
;
input
CORETSE_AHBOlo
;
input
CORETSE_AHBioOI
;
input
CORETSE_AHBOiOI
;
input
CORETSE_AHBIiOI
;
input
CORETSE_AHBliOI
;
input
CORETSE_AHBoiOI
;
output
CORETSE_AHBilII
;
output
CORETSE_AHBO0II
;
output
CORETSE_AHBI0II
;
output
CORETSE_AHBl0II
;
output
CORETSE_AHBo0II
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBloII
;
reg
CORETSE_AHBooII
;
reg
CORETSE_AHBioII
;
reg
CORETSE_AHBOiII
;
reg
CORETSE_AHBIiII
;
reg
CORETSE_AHBliII
;
reg
CORETSE_AHBoiII
;
reg
CORETSE_AHBiiII
;
reg
CORETSE_AHBOOlI
;
reg
CORETSE_AHBIOlI
;
always
@
(
posedge
CORETSE_AHBOOo
)
begin
CORETSE_AHBloII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi0
|
CORETSE_AHBioOI
;
end
always
@
(
posedge
CORETSE_AHBOOo
)
begin
CORETSE_AHBooII
<=
#
CORETSE_AHBIoII
CORETSE_AHBloII
;
end
assign
CORETSE_AHBilII
=
CORETSE_AHBoo1
?
CORETSE_AHBIi0
:
(
(
CORETSE_AHBIi0
|
CORETSE_AHBioOI
)
|
CORETSE_AHBooII
)
;
always
@
(
posedge
CORETSE_AHBOlo
)
begin
CORETSE_AHBIiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi0
|
CORETSE_AHBIiOI
;
end
always
@
(
posedge
CORETSE_AHBOlo
)
begin
CORETSE_AHBliII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIiII
;
end
assign
CORETSE_AHBI0II
=
CORETSE_AHBoo1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIiOI
|
CORETSE_AHBliII
)
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBioII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi0
|
CORETSE_AHBOiOI
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBOiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBioII
;
end
assign
CORETSE_AHBO0II
=
CORETSE_AHBoo1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBOiOI
|
CORETSE_AHBOiII
)
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBoiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi0
|
CORETSE_AHBliOI
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBiiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiII
;
end
assign
CORETSE_AHBl0II
=
CORETSE_AHBoo1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBliOI
|
CORETSE_AHBiiII
)
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBOOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi0
|
CORETSE_AHBoiOI
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBIOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOlI
;
end
assign
CORETSE_AHBo0II
=
CORETSE_AHBoo1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBoiOI
|
CORETSE_AHBIOlI
)
;
endmodule
