// REVISION    : $Revision: 1.11 $
//         Mentor Graphics Corporation Proprietary and Confidential
//         Copyright Mentor Graphics Corporation and Licensors 2004
`include "include.v"
module
decoder
(
CORETSE_AHBioOl
,
CORETSE_AHBOiOl
,
CORETSE_AHBIiOl
,
CORETSE_AHBliOl
,
CORETSE_AHBoiOl
,
CORETSE_AHBiiOl
,
CORETSE_AHBOOIl
,
CORETSE_AHBIOIl
,
CORETSE_AHBlOIl
,
CORETSE_AHBoOIl
,
CORETSE_AHBiOIl
,
CORETSE_AHBOIIl
,
CORETSE_AHBIIIl
,
CORETSE_AHBlIIl
,
CORETSE_AHBoIIl
,
CORETSE_AHBiIIl
,
CORETSE_AHBOlIl
,
CORETSE_AHBIlIl
,
CORETSE_AHBllIl
,
CORETSE_AHBolIl
,
CORETSE_AHBilIl
,
CORETSE_AHBO0Il
,
CORETSE_AHBI0Il
)
;
input
[
7
:
3
]
CORETSE_AHBOiOl
;
input
CORETSE_AHBioOl
;
output
[
31
:
0
]
CORETSE_AHBIiOl
;
output
CORETSE_AHBliOl
;
output
CORETSE_AHBoiOl
;
input
[
31
:
0
]
CORETSE_AHBiiOl
;
input
CORETSE_AHBOOIl
;
output
CORETSE_AHBIOIl
;
input
[
31
:
0
]
CORETSE_AHBlOIl
;
input
CORETSE_AHBoOIl
;
output
CORETSE_AHBiOIl
;
input
[
31
:
0
]
CORETSE_AHBOIIl
;
input
CORETSE_AHBIIIl
;
input
CORETSE_AHBlIIl
;
output
CORETSE_AHBoIIl
;
input
[
31
:
0
]
CORETSE_AHBiIIl
;
input
CORETSE_AHBOlIl
;
output
CORETSE_AHBIlIl
;
output
CORETSE_AHBilIl
;
input
CORETSE_AHBolIl
;
input
[
31
:
0
]
CORETSE_AHBllIl
;
input
CORETSE_AHBI0Il
;
input
[
31
:
0
]
CORETSE_AHBO0Il
;
wire
CORETSE_AHBl0Il
;
assign
CORETSE_AHBl0Il
=
!
(
CORETSE_AHBOiOl
[
7
:
5
]
==
`CORETSE_AHBo0Il
&
!
CORETSE_AHBioOl
)
;
assign
CORETSE_AHBIOIl
=
!
(
!
CORETSE_AHBl0Il
&
!
CORETSE_AHBOiOl
[
4
]
&
!
CORETSE_AHBioOl
)
;
assign
CORETSE_AHBiOIl
=
!
(
!
CORETSE_AHBl0Il
&
CORETSE_AHBOiOl
[
4
]
&
!
CORETSE_AHBioOl
)
;
assign
CORETSE_AHBoiOl
=
!
(
(
CORETSE_AHBOiOl
[
7
:
5
]
==
3
'b
000
)
&
!
CORETSE_AHBioOl
)
;
assign
CORETSE_AHBoIIl
=
!
(
CORETSE_AHBOiOl
[
7
:
5
]
==
`CORETSE_AHBi0Il
&
!
CORETSE_AHBioOl
)
;
assign
CORETSE_AHBilIl
=
!
(
CORETSE_AHBOiOl
[
7
:
3
]
==
`CORETSE_AHBO1Il
)
;
assign
CORETSE_AHBIlIl
=
!
(
CORETSE_AHBOiOl
[
7
:
3
]
==
`CORETSE_AHBI1Il
&
!
CORETSE_AHBioOl
)
;
assign
CORETSE_AHBIiOl
=
(
{
32
{
!
CORETSE_AHBIOIl
}
}
&
CORETSE_AHBlOIl
)
|
(
{
32
{
!
CORETSE_AHBiOIl
}
}
&
CORETSE_AHBOIIl
)
|
(
{
32
{
!
CORETSE_AHBoiOl
|
!
CORETSE_AHBlIIl
}
}
&
CORETSE_AHBiiOl
)
|
(
{
32
{
!
CORETSE_AHBoIIl
}
}
&
CORETSE_AHBiIIl
)
|
(
{
32
{
!
CORETSE_AHBIlIl
}
}
&
CORETSE_AHBllIl
)
|
(
{
32
{
!
CORETSE_AHBilIl
}
}
&
CORETSE_AHBO0Il
)
;
assign
CORETSE_AHBliOl
=
(
!
CORETSE_AHBIOIl
&
CORETSE_AHBoOIl
)
|
(
!
CORETSE_AHBiOIl
&
CORETSE_AHBIIIl
)
|
(
(
!
CORETSE_AHBoiOl
|
!
CORETSE_AHBlIIl
)
&
CORETSE_AHBOOIl
)
|
(
!
CORETSE_AHBoIIl
&
CORETSE_AHBOlIl
)
|
(
!
CORETSE_AHBIlIl
&
CORETSE_AHBolIl
)
|
(
!
CORETSE_AHBilIl
&
CORETSE_AHBI0Il
)
;
endmodule
