// REVISION    : $Revision: 1.1 $
//              Mentor Proprietary and Confidential
//              Copyright (c) 2000, Mentor Intellectual Property Development
`timescale 1ns/1ns
module
pemstat_sadd
(
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
,
CORETSE_AHBi10i
,
CORETSE_AHBOo0i
,
CORETSE_AHBoIIi
,
CORETSE_AHBl1li
,
CORETSE_AHBiIIi
,
CORETSE_AHBlIIi
,
CORETSE_AHBIo0i
,
CORETSE_AHBoOIi
)
;
input
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
;
input
CORETSE_AHBi10i
;
input
[
3
:
0
]
CORETSE_AHBOo0i
;
input
CORETSE_AHBoIIi
;
input
[
30
:
0
]
CORETSE_AHBl1li
;
input
CORETSE_AHBiIIi
;
input
CORETSE_AHBlIIi
;
output
[
30
:
0
]
CORETSE_AHBIo0i
;
output
CORETSE_AHBoOIi
;
reg
[
11
:
0
]
CORETSE_AHBoo0i
;
reg
CORETSE_AHBoOIi
;
parameter
CORETSE_AHBIoII
=
1
;
wire
[
12
:
0
]
CORETSE_AHBlo0i
;
assign
CORETSE_AHBlo0i
=
CORETSE_AHBoo0i
+
{
8
'h
0
,
CORETSE_AHBOo0i
}
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBoo0i
<=
#
CORETSE_AHBIoII
12
'h
0
;
else
if
(
CORETSE_AHBoIIi
)
CORETSE_AHBoo0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1li
[
11
:
0
]
;
else
if
(
CORETSE_AHBi10i
&
CORETSE_AHBlIIi
)
CORETSE_AHBoo0i
<=
#
CORETSE_AHBIoII
{
8
'h
0
,
CORETSE_AHBOo0i
}
;
else
if
(
CORETSE_AHBi10i
)
CORETSE_AHBoo0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo0i
[
11
:
0
]
;
else
if
(
CORETSE_AHBlIIi
)
CORETSE_AHBoo0i
<=
#
CORETSE_AHBIoII
12
'h
0
;
else
CORETSE_AHBoo0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0i
;
end
assign
CORETSE_AHBIo0i
=
{
19
'h
0
,
CORETSE_AHBoo0i
[
11
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBiIIi
)
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi10i
&
CORETSE_AHBlo0i
[
12
]
)
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOIi
;
end
endmodule
