// REVISION    : $Revision: 1.1 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_cnvtxo
(
CORETSE_AHBoO10
,
CORETSE_AHBli0
,
CORETSE_AHBo11
,
CORETSE_AHBloo0
,
CORETSE_AHBooo0
,
CORETSE_AHBioo0
,
CORETSE_AHBOio0
,
CORETSE_AHBIio0
,
CORETSE_AHBIoo0
,
CORETSE_AHBI0i0
,
CORETSE_AHBo110
,
CORETSE_AHBl0i0
,
CORETSE_AHBIl1
)
;
input
CORETSE_AHBoO10
;
input
CORETSE_AHBli0
;
input
[
1
:
0
]
CORETSE_AHBo11
;
input
[
7
:
0
]
CORETSE_AHBloo0
;
input
CORETSE_AHBooo0
;
input
CORETSE_AHBioo0
;
input
CORETSE_AHBOio0
;
input
[
2
:
0
]
CORETSE_AHBIio0
;
output
[
2
:
0
]
CORETSE_AHBIoo0
;
output
[
7
:
0
]
CORETSE_AHBI0i0
;
output
CORETSE_AHBo110
;
output
CORETSE_AHBl0i0
;
output
CORETSE_AHBIl1
;
`define CORETSE_AHBIoII  \
# \
1
reg
[
2
:
0
]
CORETSE_AHBIoo0
;
reg
[
7
:
0
]
CORETSE_AHBI0i0
;
reg
CORETSE_AHBo110
;
reg
CORETSE_AHBl0i0
;
reg
[
2
:
0
]
CORETSE_AHBO0i0
;
reg
CORETSE_AHBo0i0
;
wire
CORETSE_AHBi0i0
;
reg
[
6
:
0
]
CORETSE_AHBii10
;
wire
CORETSE_AHBO1i0
;
reg
CORETSE_AHBIl1
;
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBO0i0
<=
`CORETSE_AHBIoII
3
'h
0
;
else
CORETSE_AHBO0i0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBO0i0
[
1
:
0
]
,
CORETSE_AHBOio0
}
;
end
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBo0i0
<=
`CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBO1i0
)
CORETSE_AHBo0i0
<=
`CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBO0i0
[
2
:
1
]
==
2
'b
01
)
CORETSE_AHBo0i0
<=
`CORETSE_AHBIoII
1
'b
1
;
end
assign
CORETSE_AHBi0i0
=
(
(
CORETSE_AHBO0i0
[
2
:
1
]
==
2
'b
01
)
|
CORETSE_AHBo0i0
)
&
~
CORETSE_AHBooo0
;
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
7
'd
00
;
else
if
(
(
CORETSE_AHBo11
==
2
'b
00
)
&
CORETSE_AHBO1i0
)
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
7
'd
99
;
else
if
(
(
CORETSE_AHBo11
==
2
'b
01
)
&
CORETSE_AHBO1i0
)
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
7
'd
09
;
else
if
(
CORETSE_AHBo11
==
2
'b
10
)
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
7
'd
00
;
else
CORETSE_AHBii10
<=
`CORETSE_AHBIoII
CORETSE_AHBii10
-
7
'h
1
;
end
assign
CORETSE_AHBO1i0
=
(
CORETSE_AHBii10
==
7
'h
00
)
;
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBIoo0
<=
`CORETSE_AHBIoII
3
'h
0
;
else
if
(
CORETSE_AHBO1i0
&
CORETSE_AHBi0i0
)
CORETSE_AHBIoo0
<=
`CORETSE_AHBIoII
CORETSE_AHBIio0
;
else
if
(
CORETSE_AHBO1i0
)
CORETSE_AHBIoo0
<=
`CORETSE_AHBIoII
CORETSE_AHBIoo0
+
3
'h
1
;
end
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBIl1
<=
`CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIl1
<=
`CORETSE_AHBIoII
~
CORETSE_AHBIl1
;
end
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBI0i0
<=
`CORETSE_AHBIoII
8
'h
0
;
else
CORETSE_AHBI0i0
<=
`CORETSE_AHBIoII
CORETSE_AHBloo0
;
end
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBo110
<=
`CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo110
<=
`CORETSE_AHBIoII
CORETSE_AHBooo0
;
end
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBoO10
)
begin
if
(
CORETSE_AHBoO10
)
CORETSE_AHBl0i0
<=
`CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl0i0
<=
`CORETSE_AHBIoII
CORETSE_AHBioo0
;
end
endmodule
