// VERSION     : $Revision: 1.20 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
petfn_top
#
(
parameter
CORETSE_AHBiOI
=
0
,
parameter
CORETSE_AHBlOI
=
0
)
(
CORETSE_AHBiOO1
,
CORETSE_AHBo1Oo
,
CORETSE_AHBol
,
CORETSE_AHBll
,
CORETSE_AHBiio
,
CORETSE_AHBiOi
,
CORETSE_AHBIIi
,
CORETSE_AHBOIi
,
CORETSE_AHBoOo1
,
CORETSE_AHBilIo
,
CORETSE_AHBoo01
,
CORETSE_AHBIOOo
,
CORETSE_AHBio01
,
CORETSE_AHBi0i1
,
CORETSE_AHBlOi
,
CORETSE_AHBOOi
,
CORETSE_AHBoo11
,
CORETSE_AHBIOi
,
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
,
CORETSE_AHBIoOo
,
CORETSE_AHBlii1
,
CORETSE_AHBI1i1
,
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
,
CORETSE_AHBi1i1
,
CORETSE_AHBOoi1
,
CORETSE_AHBoii1
,
CORETSE_AHBiii1
,
CORETSE_AHBlli1
,
CORETSE_AHBIoi1
,
CORETSE_AHBiIi
,
CORETSE_AHBioi1
,
CORETSE_AHBloOo
,
CORETSE_AHBIio1
,
CORETSE_AHBlOOo
,
CORETSE_AHBloi1
,
CORETSE_AHBlOi1
,
CORETSE_AHBI0Io
,
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
,
CORETSE_AHBI0o
,
CORETSE_AHBI0o1
,
CORETSE_AHBl0o1
,
CORETSE_AHBi0o1
,
CORETSE_AHBOoo1
,
CORETSE_AHBIoo1
,
CORETSE_AHBloo1
,
CORETSE_AHBooo1
,
CORETSE_AHBioo1
,
CORETSE_AHBOio1
,
CORETSE_AHBIOo1
,
CORETSE_AHBlOo1
,
CORETSE_AHBoOi1
,
CORETSE_AHBoI
,
CORETSE_AHBII
,
CORETSE_AHBOl
)
;
input
CORETSE_AHBiOO1
,
CORETSE_AHBo1Oo
;
input
CORETSE_AHBol
,
CORETSE_AHBll
;
input
[
7
:
0
]
CORETSE_AHBiio
;
input
CORETSE_AHBiOi
,
CORETSE_AHBIIi
,
CORETSE_AHBOIi
;
input
CORETSE_AHBoOo1
,
CORETSE_AHBilIo
;
input
[
1
:
0
]
CORETSE_AHBoo01
;
input
CORETSE_AHBIOOo
,
CORETSE_AHBio01
,
CORETSE_AHBi0i1
;
input
CORETSE_AHBlOi
,
CORETSE_AHBOOi
,
CORETSE_AHBoo11
,
CORETSE_AHBIOi
;
input
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
,
CORETSE_AHBIoOo
;
input
[
3
:
0
]
CORETSE_AHBlii1
;
input
[
6
:
0
]
CORETSE_AHBI1i1
,
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
;
input
[
9
:
0
]
CORETSE_AHBi1i1
;
input
[
3
:
0
]
CORETSE_AHBOoi1
,
CORETSE_AHBoii1
;
input
CORETSE_AHBlli1
,
CORETSE_AHBloi1
;
input
CORETSE_AHBiii1
,
CORETSE_AHBIoi1
,
CORETSE_AHBiIi
,
CORETSE_AHBioi1
;
input
[
15
:
0
]
CORETSE_AHBloOo
;
input
CORETSE_AHBIio1
,
CORETSE_AHBlOOo
;
output
CORETSE_AHBlOi1
;
output
CORETSE_AHBI0Io
;
output
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
;
output
CORETSE_AHBI0o
;
output
CORETSE_AHBIOo1
;
output
[
51
:
0
]
CORETSE_AHBlOo1
;
output
CORETSE_AHBoOi1
;
output
CORETSE_AHBoI
;
output
[
7
:
0
]
CORETSE_AHBII
;
output
CORETSE_AHBOl
;
output
CORETSE_AHBI0o1
;
output
[
7
:
0
]
CORETSE_AHBl0o1
;
output
CORETSE_AHBi0o1
;
input
CORETSE_AHBOoo1
;
input
CORETSE_AHBIoo1
;
input
[
15
:
0
]
CORETSE_AHBloo1
;
input
CORETSE_AHBooo1
;
input
CORETSE_AHBOio1
;
input
[
79
:
0
]
CORETSE_AHBioo1
;
reg
CORETSE_AHBlOi1
;
reg
CORETSE_AHBI0Io
;
reg
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
;
reg
CORETSE_AHBI0o
;
reg
CORETSE_AHBIOo1
;
reg
[
51
:
0
]
CORETSE_AHBlOo1
;
reg
CORETSE_AHBoOi1
;
reg
CORETSE_AHBoI
;
reg
CORETSE_AHBi01II
;
reg
CORETSE_AHBO11II
;
wire
CORETSE_AHBI11II
;
reg
[
7
:
0
]
CORETSE_AHBII
;
reg
CORETSE_AHBOl
;
reg
CORETSE_AHBl11II
;
reg
CORETSE_AHBo11II
;
wire
CORETSE_AHBi11II
;
reg
CORETSE_AHBOo1II
;
wire
CORETSE_AHBIo1II
;
wire
CORETSE_AHBlo1II
;
wire
CORETSE_AHBoo1II
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBio1II
,
CORETSE_AHBOi1II
;
reg
CORETSE_AHBIi1II
,
CORETSE_AHBli1II
;
wire
CORETSE_AHBOilII
;
reg
CORETSE_AHBI1lOI
,
CORETSE_AHBo1lOI
;
reg
CORETSE_AHBoi1II
,
CORETSE_AHBii1II
;
wire
CORETSE_AHBOOoII
;
wire
CORETSE_AHBIOoII
;
reg
CORETSE_AHBlOoII
;
wire
CORETSE_AHBoOoII
,
CORETSE_AHBiOoII
,
CORETSE_AHBOIoII
;
reg
CORETSE_AHBIIoII
,
CORETSE_AHBlIoII
,
CORETSE_AHBO1i1
;
wire
CORETSE_AHBoIoII
;
reg
CORETSE_AHBiIoII
;
wire
CORETSE_AHBOloII
;
reg
CORETSE_AHBIloII
;
wire
CORETSE_AHBlolOI
;
reg
CORETSE_AHBoilOI
;
wire
CORETSE_AHBoolOI
;
reg
CORETSE_AHBiilOI
;
wire
CORETSE_AHBiolOI
;
reg
CORETSE_AHBOO0OI
;
wire
CORETSE_AHBlloII
,
CORETSE_AHBoloII
;
reg
CORETSE_AHBiloII
,
CORETSE_AHBO0oII
;
wire
CORETSE_AHBI0oII
;
reg
CORETSE_AHBl0oII
;
wire
CORETSE_AHBo0oII
;
reg
CORETSE_AHBi0oII
;
wire
CORETSE_AHBO1oII
;
reg
CORETSE_AHBI1oII
;
wire
CORETSE_AHBl1oII
;
reg
CORETSE_AHBo1oII
;
wire
CORETSE_AHBi1oII
;
reg
CORETSE_AHBOooII
;
reg
CORETSE_AHBIooII
;
reg
CORETSE_AHBlooII
;
wire
CORETSE_AHBoooII
;
reg
CORETSE_AHBiooII
;
reg
[
3
:
0
]
CORETSE_AHBOioII
;
reg
[
15
:
0
]
CORETSE_AHBIioII
;
reg
CORETSE_AHBlioII
,
CORETSE_AHBoioII
,
CORETSE_AHBiioII
;
reg
CORETSE_AHBOOiII
,
CORETSE_AHBIOiII
;
wire
[
3
:
0
]
CORETSE_AHBlOiII
;
reg
[
3
:
0
]
CORETSE_AHBoOiII
;
reg
[
3
:
0
]
CORETSE_AHBiOiII
;
reg
[
3
:
0
]
CORETSE_AHBOIiII
;
wire
[
3
:
0
]
CORETSE_AHBIIiII
;
wire
CORETSE_AHBlIiII
;
wire
CORETSE_AHBoIiII
,
CORETSE_AHBiIiII
;
reg
CORETSE_AHBOliII
,
CORETSE_AHBIliII
,
CORETSE_AHBlliII
;
wire
[
7
:
0
]
CORETSE_AHBoliII
;
wire
CORETSE_AHBiliII
;
reg
CORETSE_AHBO0iII
;
wire
CORETSE_AHBI0iII
;
reg
CORETSE_AHBl0iII
;
wire
CORETSE_AHBo0iII
;
reg
CORETSE_AHBi0iII
;
wire
CORETSE_AHBO1iII
;
wire
CORETSE_AHBI1iII
;
reg
CORETSE_AHBl1iII
,
CORETSE_AHBo1iII
;
reg
CORETSE_AHBi1iII
;
wire
CORETSE_AHBOoiII
,
CORETSE_AHBIoiII
;
wire
[
6
:
0
]
CORETSE_AHBloiII
;
reg
[
6
:
0
]
CORETSE_AHBooiII
;
wire
[
6
:
0
]
CORETSE_AHBioiII
;
reg
[
6
:
0
]
CORETSE_AHBOiiII
;
wire
CORETSE_AHBIiiII
,
CORETSE_AHBliiII
;
wire
[
3
:
0
]
CORETSE_AHBoiiII
;
reg
[
3
:
0
]
CORETSE_AHBiiiII
;
wire
CORETSE_AHBOOOlI
,
CORETSE_AHBIOOlI
;
wire
[
15
:
0
]
CORETSE_AHBlOOlI
;
reg
[
15
:
0
]
CORETSE_AHBoOOlI
;
wire
CORETSE_AHBil0OI
,
CORETSE_AHBO00OI
,
CORETSE_AHBI00OI
;
wire
CORETSE_AHBl00OI
,
CORETSE_AHBo00OI
,
CORETSE_AHBO10OI
;
wire
CORETSE_AHBl10OI
,
CORETSE_AHBo1oOI
,
CORETSE_AHBo10OI
;
wire
CORETSE_AHBOo0OI
,
CORETSE_AHBiOOlI
;
wire
CORETSE_AHBOIOlI
;
wire
CORETSE_AHBIIOlI
;
wire
CORETSE_AHBlIOlI
,
CORETSE_AHBoIOlI
;
wire
[
15
:
0
]
CORETSE_AHBiIOlI
;
reg
[
15
:
0
]
CORETSE_AHBOlOlI
;
wire
CORETSE_AHBIlOlI
;
reg
CORETSE_AHBllOlI
;
wire
CORETSE_AHBolOlI
,
CORETSE_AHBilOlI
;
wire
[
3
:
0
]
CORETSE_AHBO0OlI
;
reg
[
3
:
0
]
CORETSE_AHBI0OlI
;
wire
CORETSE_AHBl0OlI
;
wire
[
11
:
1
]
CORETSE_AHBo0OlI
;
reg
[
11
:
1
]
CORETSE_AHBi0OlI
;
wire
CORETSE_AHBO1OlI
;
wire
[
9
:
0
]
CORETSE_AHBI1OlI
;
reg
[
9
:
0
]
CORETSE_AHBl1OlI
;
wire
CORETSE_AHBo1OlI
,
CORETSE_AHBi1OlI
;
wire
[
10
:
1
]
CORETSE_AHBOoOlI
;
wire
CORETSE_AHBIli1
,
CORETSE_AHBIoOlI
;
wire
[
8
:
0
]
CORETSE_AHBOIOII
;
reg
[
8
:
0
]
CORETSE_AHBIIOII
;
wire
CORETSE_AHBloOlI
,
CORETSE_AHBooOlI
;
wire
[
9
:
0
]
CORETSE_AHBioOlI
;
reg
[
9
:
0
]
CORETSE_AHBOiOlI
;
reg
CORETSE_AHBIiOlI
;
wire
CORETSE_AHBliOlI
,
CORETSE_AHBoiOlI
,
CORETSE_AHBiiOlI
,
CORETSE_AHBOOIlI
;
reg
CORETSE_AHBIOIlI
;
wire
CORETSE_AHBillII
;
wire
CORETSE_AHBlOIlI
;
reg
CORETSE_AHBO0lII
;
wire
[
7
:
0
]
CORETSE_AHBoOIlI
;
reg
[
7
:
0
]
CORETSE_AHBiOIlI
;
wire
[
7
:
0
]
CORETSE_AHBOIIlI
;
wire
[
7
:
0
]
CORETSE_AHBIIIlI
;
reg
[
7
:
0
]
CORETSE_AHBlIIlI
;
wire
[
7
:
0
]
CORETSE_AHBoIIlI
;
reg
[
7
:
0
]
CORETSE_AHBiIIlI
;
reg
[
7
:
0
]
CORETSE_AHBOlIlI
;
wire
[
7
:
0
]
CORETSE_AHBIlIlI
;
wire
[
7
:
0
]
CORETSE_AHBllIlI
;
wire
CORETSE_AHBI11OI
,
CORETSE_AHBl11OI
,
CORETSE_AHBo11OI
;
reg
CORETSE_AHBil1o
,
CORETSE_AHBolIlI
,
CORETSE_AHBilIlI
,
CORETSE_AHBol1o
,
CORETSE_AHBO0IlI
,
CORETSE_AHBI0IlI
,
CORETSE_AHBO01o
,
CORETSE_AHBl0IlI
,
CORETSE_AHBo0IlI
;
wire
CORETSE_AHBi0IlI
,
CORETSE_AHBO1IlI
,
CORETSE_AHBI1IlI
;
wire
[
31
:
0
]
CORETSE_AHBl01o
;
wire
CORETSE_AHBo01o
;
wire
[
7
:
0
]
CORETSE_AHBl1IlI
,
CORETSE_AHBo1IlI
,
CORETSE_AHBi1IlI
,
CORETSE_AHBOoIlI
;
wire
CORETSE_AHBIoIlI
;
wire
[
7
:
0
]
CORETSE_AHBloIlI
;
wire
[
7
:
0
]
CORETSE_AHBooIlI
;
wire
CORETSE_AHBioIlI
;
wire
CORETSE_AHBii0OI
,
CORETSE_AHBOiIlI
;
wire
CORETSE_AHBIiIlI
,
CORETSE_AHBliIlI
,
CORETSE_AHBoiIlI
,
CORETSE_AHBiiIlI
;
reg
CORETSE_AHBOOllI
,
CORETSE_AHBIOllI
;
reg
CORETSE_AHBlOllI
,
CORETSE_AHBoOllI
,
CORETSE_AHBiOllI
,
CORETSE_AHBOIllI
;
wire
CORETSE_AHBIIllI
,
CORETSE_AHBlIllI
;
reg
CORETSE_AHBoIllI
,
CORETSE_AHBiIllI
,
CORETSE_AHBOlllI
;
wire
CORETSE_AHBIlllI
;
reg
CORETSE_AHBllllI
;
wire
CORETSE_AHBolllI
;
reg
CORETSE_AHBilllI
;
wire
CORETSE_AHBO0llI
;
reg
CORETSE_AHBI0llI
;
wire
CORETSE_AHBIo1OI
,
CORETSE_AHBlo1OI
;
reg
CORETSE_AHBOl00
,
CORETSE_AHBiI00
;
wire
CORETSE_AHBoo1OI
,
CORETSE_AHBio1OI
;
wire
[
15
:
0
]
CORETSE_AHBOi1OI
;
reg
[
15
:
0
]
CORETSE_AHBIi1OI
;
wire
CORETSE_AHBli1OI
,
CORETSE_AHBoi1OI
,
CORETSE_AHBl0llI
;
wire
CORETSE_AHBii1OI
;
reg
CORETSE_AHBOOoOI
;
wire
CORETSE_AHBo0llI
;
reg
CORETSE_AHBi0llI
;
wire
[
15
:
0
]
CORETSE_AHBiOoOI
;
wire
CORETSE_AHBOIoOI
,
CORETSE_AHBO1llI
;
reg
CORETSE_AHBIIoOI
;
wire
CORETSE_AHBI1llI
,
CORETSE_AHBl1llI
;
reg
CORETSE_AHBo1llI
,
CORETSE_AHBi1llI
;
wire
CORETSE_AHBOollI
;
wire
[
51
:
0
]
CORETSE_AHBIollI
;
reg
[
9
:
0
]
CORETSE_AHBlollI
;
assign
CORETSE_AHBI0o1
=
CORETSE_AHBo1llI
;
assign
CORETSE_AHBi0o1
=
CORETSE_AHBOO0OI
;
assign
CORETSE_AHBl0o1
=
CORETSE_AHBoOIlI
;
assign
CORETSE_AHBOIIlI
=
CORETSE_AHBiOIlI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIi1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIi1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOOo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBli1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBli1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi1II
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlOi1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlOi1
<=
#
CORETSE_AHBIoII
~
CORETSE_AHBO0lII
&
CORETSE_AHBli1II
|
CORETSE_AHBO0lII
&
CORETSE_AHBlOi1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBI1lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI1lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBo1lOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo1lOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1lOI
&
~
CORETSE_AHBio01
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBoi1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoi1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBll
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBii1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBii1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBoi1II
;
end
assign
CORETSE_AHBOOoII
=
CORETSE_AHBiilOI
|
CORETSE_AHBOO0OI
|
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
|
CORETSE_AHBl0oII
|
CORETSE_AHBI1oII
;
assign
CORETSE_AHBIOoII
=
CORETSE_AHBOOoII
&
(
~
CORETSE_AHBlOoII
&
CORETSE_AHBii1II
&
~
CORETSE_AHBio01
|
CORETSE_AHBlOoII
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlOoII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlOoII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOoII
;
end
assign
CORETSE_AHBoOoII
=
~
CORETSE_AHBIIoII
&
CORETSE_AHBiOi
&
CORETSE_AHBolo
&
(
CORETSE_AHBl0i1
|
CORETSE_AHBIOi
&
CORETSE_AHBlOi
|
CORETSE_AHBoOo1
)
|
CORETSE_AHBIIoII
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIIoII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIIoII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOoII
;
end
assign
CORETSE_AHBiOoII
=
CORETSE_AHBiOi
&
CORETSE_AHBolo
&
(
CORETSE_AHBl0i1
|
CORETSE_AHBo0i1
|
CORETSE_AHBIOi
&
(
CORETSE_AHBlOi
|
CORETSE_AHBOOi
)
|
CORETSE_AHBoOo1
)
|
~
(
CORETSE_AHBiOi
&
CORETSE_AHBolo
)
&
CORETSE_AHBlIoII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlIoII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBlIoII
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOoII
;
end
assign
CORETSE_AHBOIoII
=
CORETSE_AHBiOi
&
CORETSE_AHBolo
&
(
CORETSE_AHBIoOo
|
CORETSE_AHBIOi
&
CORETSE_AHBoo11
)
|
~
(
CORETSE_AHBiOi
&
CORETSE_AHBolo
)
&
CORETSE_AHBO1i1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBO1i1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO1i1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIoII
;
end
assign
CORETSE_AHBoIoII
=
CORETSE_AHBiIoII
&
(
CORETSE_AHBo1lOI
|
~
CORETSE_AHBlOi1
)
|
CORETSE_AHBIloII
&
CORETSE_AHBo1lOI
&
CORETSE_AHBooiII
[
6
:
0
]
>
CORETSE_AHBOiiII
[
6
:
0
]
|
CORETSE_AHBoilOI
&
CORETSE_AHBo1lOI
&
~
CORETSE_AHBiOi
|
CORETSE_AHBiilOI
&
(
~
CORETSE_AHBl1iII
&
CORETSE_AHBo1iII
|
CORETSE_AHBl1iII
&
(
&
CORETSE_AHBOlOlI
[
11
:
0
]
)
)
|
CORETSE_AHBiloII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
&
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBO0oII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
&
~
CORETSE_AHBOliII
|
CORETSE_AHBOliII
&
CORETSE_AHBlIiII
&
(
CORETSE_AHBo1OlI
|
~
CORETSE_AHBllOlI
|
CORETSE_AHBl0OlI
|
CORETSE_AHBO1iII
)
|
CORETSE_AHBO0iII
&
(
CORETSE_AHBi1OlI
|
CORETSE_AHBIIi
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiIoII
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiIoII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIoII
;
end
assign
CORETSE_AHBOloII
=
CORETSE_AHBiIoII
&
~
CORETSE_AHBo1lOI
&
CORETSE_AHBlOi1
|
CORETSE_AHBIloII
&
(
CORETSE_AHBl0iII
&
|
CORETSE_AHBooiII
[
6
:
0
]
|
~
CORETSE_AHBl0iII
&
|
CORETSE_AHBooiII
[
6
:
0
]
)
&
~
(
CORETSE_AHBo1lOI
&
CORETSE_AHBooiII
[
6
:
0
]
>
CORETSE_AHBOiiII
[
6
:
0
]
)
&
~
CORETSE_AHBl1iII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIloII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIloII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOloII
;
end
assign
CORETSE_AHBlolOI
=
CORETSE_AHBIloII
&
(
CORETSE_AHBl0iII
&
~|
CORETSE_AHBooiII
[
6
:
0
]
|
~
CORETSE_AHBl0iII
&
~|
CORETSE_AHBooiII
[
6
:
0
]
)
|
CORETSE_AHBoilOI
&
~
(
CORETSE_AHBiOi
|
CORETSE_AHBo1lOI
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBoilOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoilOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlolOI
;
end
assign
CORETSE_AHBoolOI
=
CORETSE_AHBoilOI
&
CORETSE_AHBiOi
|
CORETSE_AHBl1iII
|
CORETSE_AHBiilOI
&
|
CORETSE_AHBiiiII
[
3
:
0
]
&
~
(
~
CORETSE_AHBl1iII
&
CORETSE_AHBo1iII
|
CORETSE_AHBl1iII
&
(
&
CORETSE_AHBOlOlI
[
11
:
0
]
)
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiilOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiilOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoolOI
;
end
assign
CORETSE_AHBiolOI
=
CORETSE_AHBiilOI
&
CORETSE_AHBiiiII
[
3
:
0
]
==
4
'h
1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOO0OI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOO0OI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiolOI
;
end
assign
CORETSE_AHBlloII
=
CORETSE_AHBiilOI
&
~
CORETSE_AHBlOoII
&
~|
CORETSE_AHBiiiII
[
3
:
0
]
|
CORETSE_AHBO0oII
&
~
CORETSE_AHBlOoII
&
~
CORETSE_AHBOIi
&
~
CORETSE_AHBOOllI
&
~
CORETSE_AHBIOllI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiloII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiloII
<=
#
CORETSE_AHBIoII
CORETSE_AHBlloII
;
end
assign
CORETSE_AHBoloII
=
CORETSE_AHBiloII
&
~
CORETSE_AHBlOoII
&
~
CORETSE_AHBIIi
&
~
CORETSE_AHBOOllI
&
~
CORETSE_AHBIOllI
&
~
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBiloII
&
~
CORETSE_AHBlOoII
&
~
CORETSE_AHBOIi
&
~
CORETSE_AHBIIi
&
~
CORETSE_AHBOOllI
&
~
CORETSE_AHBIOllI
&
CORETSE_AHBoo01
[
1
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBO0oII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO0oII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoloII
;
end
assign
CORETSE_AHBI0oII
=
(
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
)
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
CORETSE_AHBIIoII
&
CORETSE_AHBoOOlI
[
15
:
0
]
<
16
'h
003b
|
CORETSE_AHBl0oII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBoOOlI
[
15
:
0
]
<
16
'h
003b
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBl0oII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBl0oII
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0oII
;
end
assign
CORETSE_AHBo0oII
=
~
CORETSE_AHBO0oII
&
~
CORETSE_AHBl0oII
|
~
CORETSE_AHBi0oII
&
CORETSE_AHBl0oII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBi0oII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi0oII
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0oII
;
end
assign
CORETSE_AHBO1oII
=
(
CORETSE_AHBiloII
&
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBO0oII
)
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
(
CORETSE_AHBlIoII
&
~
CORETSE_AHBIIoII
|
CORETSE_AHBIIoII
&
CORETSE_AHBoOOlI
[
15
:
0
]
>=
16
'h
003b
)
|
CORETSE_AHBl0oII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
003b
|
CORETSE_AHBI1oII
&
~
CORETSE_AHBlIiII
|
CORETSE_AHBoIiII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBI1oII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBI1oII
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1oII
;
end
assign
CORETSE_AHBl1oII
=
~
CORETSE_AHBo1oII
&
CORETSE_AHBI1oII
|
CORETSE_AHBo1oII
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBo1oII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBo1oII
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1oII
;
end
assign
CORETSE_AHBi1oII
=
CORETSE_AHBoo01
!=
2
'h
0
&
~
CORETSE_AHBO0oII
&
~
CORETSE_AHBI1oII
|
CORETSE_AHBoo01
==
2
'h
0
&
~
CORETSE_AHBiloII
&
~
CORETSE_AHBI1oII
|
~
CORETSE_AHBOooII
&
CORETSE_AHBI1oII
|
CORETSE_AHBl1iII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBOooII
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBIooII
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBlooII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBOooII
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1oII
;
CORETSE_AHBIooII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOooII
;
CORETSE_AHBlooII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoooII
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBiooII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBiooII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIooII
;
end
end
assign
CORETSE_AHBoooII
=
CORETSE_AHBiooII
;
assign
CORETSE_AHBlOiII
[
3
:
0
]
=
{
4
{
CORETSE_AHBoo01
[
1
]
|
~
CORETSE_AHBOooII
}
}
&
{
CORETSE_AHBI1oII
&
~|
CORETSE_AHBoOiII
[
3
:
0
]
,
CORETSE_AHBoOiII
[
3
:
1
]
}
|
{
4
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOooII
}
}
&
CORETSE_AHBoOiII
[
3
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBoOiII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
4
'b
0000
;
CORETSE_AHBiOiII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
4
'b
0000
;
CORETSE_AHBOIiII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
4
'b
0000
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBoOiII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOiII
[
3
:
0
]
;
CORETSE_AHBiOiII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOiII
[
3
:
0
]
;
CORETSE_AHBOIiII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIiII
[
3
:
0
]
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBOioII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
4
'b
0000
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBOioII
[
3
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiII
[
3
:
0
]
;
end
end
assign
CORETSE_AHBIIiII
=
CORETSE_AHBOioII
;
assign
CORETSE_AHBlIiII
=
(
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBoOiII
[
1
]
|
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBoOiII
[
0
]
)
;
assign
CORETSE_AHBoIiII
=
CORETSE_AHBiilOI
&
CORETSE_AHBlOoII
&
~|
CORETSE_AHBiiiII
[
3
:
0
]
|
CORETSE_AHBiloII
&
CORETSE_AHBlOoII
|
CORETSE_AHBO0oII
&
CORETSE_AHBlOoII
|
CORETSE_AHBl0oII
&
CORETSE_AHBlOoII
|
CORETSE_AHBI1oII
&
CORETSE_AHBlOoII
&
~|
CORETSE_AHBoOiII
[
3
:
0
]
|
CORETSE_AHBii0OI
|
CORETSE_AHBOiIlI
;
assign
CORETSE_AHBiIiII
=
CORETSE_AHBoIiII
|
CORETSE_AHBOliII
&
CORETSE_AHBI1oII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBOliII
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBIliII
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBlliII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBOliII
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIiII
;
CORETSE_AHBIliII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOliII
;
CORETSE_AHBlliII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIliII
;
end
end
assign
CORETSE_AHBoliII
=
{
8
{
CORETSE_AHBlliII
}
}
&
8
'h
FF
;
assign
CORETSE_AHBiliII
=
CORETSE_AHBOliII
&
CORETSE_AHBllOlI
&
~
CORETSE_AHBo1OlI
&
~
CORETSE_AHBl0OlI
&
~
CORETSE_AHBO1iII
&
CORETSE_AHBlIiII
|
CORETSE_AHBO0iII
&
~
(
CORETSE_AHBi1OlI
|
CORETSE_AHBIIi
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBO0iII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO0iII
<=
#
CORETSE_AHBIoII
CORETSE_AHBiliII
;
end
assign
CORETSE_AHBI0iII
=
CORETSE_AHBio01
|
~
CORETSE_AHBl0iII
&
CORETSE_AHBiilOI
|
CORETSE_AHBl0iII
&
~
CORETSE_AHBiIoII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBl0iII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBl0iII
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0iII
;
end
assign
CORETSE_AHBo0iII
=
~
CORETSE_AHBi0iII
&
CORETSE_AHBiIoII
&
CORETSE_AHBo1lOI
&
CORETSE_AHBiOi
&
~
CORETSE_AHBO0lII
|
CORETSE_AHBi0iII
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBi0iII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi0iII
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0iII
;
end
assign
CORETSE_AHBO1iII
=
CORETSE_AHBIoi1
|
CORETSE_AHBiIi
&
CORETSE_AHBioi1
;
assign
CORETSE_AHBIlllI
=
CORETSE_AHBiIi
&
~
CORETSE_AHBllllI
|
CORETSE_AHBllllI
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBllllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBllllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIlllI
;
end
assign
CORETSE_AHBI1iII
=
~
CORETSE_AHBl1iII
&
CORETSE_AHBoilOI
&
CORETSE_AHBiIi
&
~
CORETSE_AHBiOi
&
~
CORETSE_AHBO0lII
|
~
CORETSE_AHBl1iII
&
CORETSE_AHBIloII
&
CORETSE_AHBiIi
&
~
CORETSE_AHBiOi
&
CORETSE_AHBooiII
[
6
:
0
]
<=
7
'h
0a
|
CORETSE_AHBl1iII
&
CORETSE_AHBiIi
&
~
CORETSE_AHBiOi
&
~&
CORETSE_AHBOlOlI
[
11
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBl1iII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBl1iII
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1iII
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBo1iII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBo1iII
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1iII
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBi1iII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi1iII
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1iII
&
~
CORETSE_AHBi1iII
;
end
assign
CORETSE_AHBOoiII
=
CORETSE_AHBiIoII
&
~
CORETSE_AHBo1lOI
;
assign
CORETSE_AHBIoiII
=
CORETSE_AHBIloII
;
assign
CORETSE_AHBloiII
[
6
:
0
]
=
{
7
{
CORETSE_AHBOoiII
&
CORETSE_AHBl0iII
&
CORETSE_AHBoo01
==
2
'b
01
}
}
&
CORETSE_AHBI1i1
[
6
:
2
]
-
2
'h
3
|
{
7
{
CORETSE_AHBOoiII
&
CORETSE_AHBl0iII
&
CORETSE_AHBoo01
==
2
'b
10
}
}
&
CORETSE_AHBI1i1
[
6
:
3
]
-
2
'h
3
|
{
7
{
CORETSE_AHBOoiII
&
~
CORETSE_AHBl0iII
&
CORETSE_AHBoo01
==
2
'b
01
}
}
&
CORETSE_AHBo1i1
[
6
:
2
]
-
3
'h
7
|
{
7
{
CORETSE_AHBOoiII
&
~
CORETSE_AHBl0iII
&
CORETSE_AHBoo01
==
2
'b
10
}
}
&
CORETSE_AHBo1i1
[
6
:
3
]
-
3
'h
7
|
{
7
{
~
CORETSE_AHBOoiII
&
CORETSE_AHBIoiII
}
}
&
CORETSE_AHBooiII
[
6
:
0
]
-
1
'b
1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBooiII
<=
#
CORETSE_AHBIoII
7
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBooiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBloiII
[
6
:
0
]
;
end
assign
CORETSE_AHBioiII
[
6
:
0
]
=
{
7
{
CORETSE_AHBoo01
==
2
'b
01
}
}
&
CORETSE_AHBl1i1
[
6
:
2
]
|
{
7
{
CORETSE_AHBoo01
==
2
'b
10
}
}
&
CORETSE_AHBl1i1
[
6
:
3
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOiiII
<=
#
CORETSE_AHBIoII
7
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOiiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBioiII
[
6
:
0
]
;
end
assign
CORETSE_AHBIiiII
=
~
CORETSE_AHBiilOI
|
CORETSE_AHBl1iII
;
assign
CORETSE_AHBliiII
=
CORETSE_AHBiilOI
;
assign
CORETSE_AHBoiiII
[
3
:
0
]
=
{
4
{
CORETSE_AHBIiiII
&
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBlii1
[
3
:
0
]
|
{
4
{
CORETSE_AHBIiiII
&
~
CORETSE_AHBoo01
[
1
]
}
}
&
{
CORETSE_AHBlii1
[
2
:
0
]
,
1
'b
1
}
|
{
4
{
~
CORETSE_AHBIiiII
&
CORETSE_AHBliiII
}
}
&
CORETSE_AHBiiiII
[
3
:
0
]
-
1
'b
1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiiiII
<=
#
CORETSE_AHBIoII
4
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiiiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiiII
[
3
:
0
]
;
end
assign
CORETSE_AHBOOOlI
=
CORETSE_AHBiilOI
|
CORETSE_AHBOollI
;
assign
CORETSE_AHBIOOlI
=
~
(
&
CORETSE_AHBoOOlI
[
15
:
0
]
)
&
(
CORETSE_AHBiIoII
&
CORETSE_AHBo1lOI
&
CORETSE_AHBiOi
&
~
CORETSE_AHBO0lII
|
CORETSE_AHBiloII
&
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBO0oII
|
CORETSE_AHBl0oII
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBi0oII
)
|
CORETSE_AHBI1oII
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBOooII
)
)
;
assign
CORETSE_AHBlOOlI
[
15
:
0
]
=
{
16
{
~
CORETSE_AHBOOOlI
&
CORETSE_AHBIOOlI
}
}
&
CORETSE_AHBoOOlI
[
15
:
0
]
+
1
'b
1
|
{
16
{
~
CORETSE_AHBOOOlI
&
~
CORETSE_AHBIOOlI
}
}
&
CORETSE_AHBoOOlI
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBoOOlI
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoOOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOOlI
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIioII
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIioII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOOlI
[
15
:
0
]
;
end
assign
CORETSE_AHBil0OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0001
;
assign
CORETSE_AHBO00OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0002
;
assign
CORETSE_AHBI00OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0003
;
assign
CORETSE_AHBl00OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0004
;
assign
CORETSE_AHBo00OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0005
;
assign
CORETSE_AHBO10OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0006
;
assign
CORETSE_AHBOIOlI
=
CORETSE_AHBoOOlI
[
15
:
0
]
>
16
'h
0006
;
assign
CORETSE_AHBl10OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
000d
;
assign
CORETSE_AHBo1oOI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
000e
;
assign
CORETSE_AHBo10OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
000f
;
assign
CORETSE_AHBOo0OI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0011
;
assign
CORETSE_AHBiOOlI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0012
;
assign
CORETSE_AHBIIOlI
=
CORETSE_AHBoOOlI
[
15
:
0
]
==
CORETSE_AHBloOo
[
15
:
0
]
&
~
CORETSE_AHBO1i1
;
assign
CORETSE_AHBlIOlI
=
CORETSE_AHBi1llI
;
assign
CORETSE_AHBoIOlI
=
~
(
&
CORETSE_AHBOlOlI
[
15
:
0
]
)
&
(
CORETSE_AHBiloII
&
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBO0oII
|
CORETSE_AHBl0oII
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBi0oII
)
|
CORETSE_AHBI1oII
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBOooII
)
|
CORETSE_AHBi1iII
)
;
assign
CORETSE_AHBiIOlI
[
15
:
0
]
=
{
16
{
~
CORETSE_AHBlIOlI
&
CORETSE_AHBoIOlI
}
}
&
CORETSE_AHBOlOlI
[
15
:
0
]
+
1
'b
1
|
{
16
{
~
CORETSE_AHBlIOlI
&
~
CORETSE_AHBoIOlI
}
}
&
CORETSE_AHBOlOlI
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOlOlI
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOlOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIOlI
[
15
:
0
]
;
end
assign
CORETSE_AHBIlOlI
=
~
CORETSE_AHBllOlI
&
~
CORETSE_AHBio01
&
CORETSE_AHBoilOI
&
CORETSE_AHBiOi
|
CORETSE_AHBllOlI
&
~
(
~
CORETSE_AHBlOoII
&
CORETSE_AHBoOOlI
[
5
:
0
]
==
CORETSE_AHBi1i1
[
5
:
0
]
&
(
CORETSE_AHBiloII
&
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBO0oII
|
CORETSE_AHBl0oII
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBi0oII
)
|
CORETSE_AHBI1oII
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBOooII
)
&
~
CORETSE_AHBOliII
)
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBllOlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBllOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIlOlI
;
end
assign
CORETSE_AHBilOlI
=
CORETSE_AHBO0iII
&
CORETSE_AHBi1OlI
|
CORETSE_AHBOliII
&
CORETSE_AHBllOlI
&
(
CORETSE_AHBo1OlI
|
CORETSE_AHBO1iII
)
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
;
assign
CORETSE_AHBolOlI
=
CORETSE_AHBIOo1
|
CORETSE_AHBOOllI
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
|
CORETSE_AHBIOllI
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
;
assign
CORETSE_AHBO0OlI
[
3
:
0
]
=
{
4
{
CORETSE_AHBilOlI
&
~
CORETSE_AHBolOlI
}
}
&
CORETSE_AHBI0OlI
[
3
:
0
]
+
1
'b
1
|
{
4
{
~
CORETSE_AHBilOlI
&
~
CORETSE_AHBolOlI
}
}
&
CORETSE_AHBI0OlI
[
3
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBI0OlI
<=
#
CORETSE_AHBIoII
4
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBI0OlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0OlI
[
3
:
0
]
;
end
assign
CORETSE_AHBl0OlI
=
CORETSE_AHBI0OlI
[
3
:
0
]
==
CORETSE_AHBOoi1
[
3
:
0
]
;
assign
CORETSE_AHBo0OlI
[
11
:
1
]
=
{
11
{
~
CORETSE_AHBlOOo
&
~
CORETSE_AHBlli1
}
}
&
{
CORETSE_AHBi0OlI
[
6
:
3
]
,
CORETSE_AHBi0OlI
[
2
]
^
(
CORETSE_AHBl01o
[
2
]
&
CORETSE_AHBO0oII
)
,
CORETSE_AHBi0OlI
[
1
]
|
CORETSE_AHBi0OlI
[
11
:
2
]
==
10
'h
0
,
CORETSE_AHBi0OlI
[
11
:
7
]
^
CORETSE_AHBi0OlI
[
9
:
5
]
}
|
{
11
{
~
CORETSE_AHBlOOo
&
CORETSE_AHBlli1
}
}
&
11
'h
7FF
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBi0OlI
<=
#
CORETSE_AHBIoII
11
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi0OlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0OlI
[
11
:
1
]
;
end
assign
CORETSE_AHBO1OlI
=
CORETSE_AHBOliII
&
CORETSE_AHBoOiII
[
3
]
&
CORETSE_AHBOooII
;
assign
CORETSE_AHBI1OlI
[
9
:
0
]
=
{
10
{
CORETSE_AHBO1OlI
}
}
&
{
CORETSE_AHBi0OlI
[
10
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
9
&
CORETSE_AHBOoOlI
[
10
]
,
CORETSE_AHBi0OlI
[
9
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
8
&
CORETSE_AHBOoOlI
[
9
]
,
CORETSE_AHBi0OlI
[
8
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
7
&
CORETSE_AHBOoOlI
[
8
]
,
CORETSE_AHBi0OlI
[
7
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
6
&
CORETSE_AHBOoOlI
[
7
]
,
CORETSE_AHBi0OlI
[
6
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
5
&
CORETSE_AHBOoOlI
[
6
]
,
CORETSE_AHBi0OlI
[
5
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
4
&
CORETSE_AHBOoOlI
[
5
]
,
CORETSE_AHBi0OlI
[
4
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
3
&
CORETSE_AHBOoOlI
[
4
]
,
CORETSE_AHBi0OlI
[
3
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
2
&
CORETSE_AHBOoOlI
[
3
]
,
CORETSE_AHBi0OlI
[
2
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
1
&
CORETSE_AHBOoOlI
[
2
]
,
CORETSE_AHBi0OlI
[
1
]
&
CORETSE_AHBI0OlI
[
3
:
0
]
>=
4
'h
0
&
CORETSE_AHBOoOlI
[
1
]
}
|
{
10
{
~
CORETSE_AHBO1OlI
}
}
&
CORETSE_AHBl1OlI
[
9
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBl1OlI
<=
#
CORETSE_AHBIoII
10
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBl1OlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1OlI
[
9
:
0
]
;
end
assign
CORETSE_AHBo1OlI
=
CORETSE_AHBl1OlI
[
9
:
0
]
==
10
'h
0
;
assign
CORETSE_AHBi1OlI
=
CORETSE_AHBOiOlI
[
9
:
0
]
==
CORETSE_AHBl1OlI
[
9
:
0
]
;
assign
CORETSE_AHBOoOlI
[
10
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
A
)
;
assign
CORETSE_AHBOoOlI
[
9
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
9
)
;
assign
CORETSE_AHBOoOlI
[
8
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
8
)
;
assign
CORETSE_AHBOoOlI
[
7
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
7
)
;
assign
CORETSE_AHBOoOlI
[
6
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
6
)
;
assign
CORETSE_AHBOoOlI
[
5
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
5
)
;
assign
CORETSE_AHBOoOlI
[
4
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
4
)
;
assign
CORETSE_AHBOoOlI
[
3
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
3
)
;
assign
CORETSE_AHBOoOlI
[
2
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
2
)
;
assign
CORETSE_AHBOoOlI
[
1
]
=
(
~
CORETSE_AHBiii1
|
CORETSE_AHBiii1
&
CORETSE_AHBoii1
[
3
:
0
]
>=
4
'h
1
)
;
assign
CORETSE_AHBIli1
=
CORETSE_AHBO0iII
&
(
&
CORETSE_AHBIIOII
[
8
:
0
]
)
;
assign
CORETSE_AHBIoOlI
=
CORETSE_AHBO0iII
;
assign
CORETSE_AHBOIOII
[
8
:
0
]
=
{
9
{
CORETSE_AHBIli1
&
CORETSE_AHBOiOlI
==
10
'h
0
}
}
&
(
{
~|
CORETSE_AHBoo01
[
1
:
0
]
,
~|
CORETSE_AHBoo01
[
1
:
0
]
,
CORETSE_AHBoo01
[
0
]
,
6
'b
11_1101
}
-
9
'h
18
)
|
{
9
{
CORETSE_AHBIli1
&
CORETSE_AHBOiOlI
!=
10
'h
0
}
}
&
{
~|
CORETSE_AHBoo01
[
1
:
0
]
,
~|
CORETSE_AHBoo01
[
1
:
0
]
,
CORETSE_AHBoo01
[
0
]
,
6
'b
11_1110
}
|
{
9
{
~
CORETSE_AHBIli1
&
CORETSE_AHBIoOlI
}
}
&
CORETSE_AHBIIOII
[
8
:
0
]
-
1
'b
1
|
{
9
{
~
CORETSE_AHBIli1
&
~
CORETSE_AHBIoOlI
}
}
&
9
'h
1ff
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIIOII
<=
#
CORETSE_AHBIoII
9
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIIOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIOII
[
8
:
0
]
;
end
assign
CORETSE_AHBloOlI
=
CORETSE_AHBoilOI
;
assign
CORETSE_AHBooOlI
=
CORETSE_AHBO0iII
&
~|
CORETSE_AHBIIOII
[
8
:
0
]
;
assign
CORETSE_AHBioOlI
[
9
:
0
]
=
{
10
{
CORETSE_AHBooOlI
}
}
&
CORETSE_AHBOiOlI
[
9
:
0
]
+
1
'b
1
|
{
10
{
~
CORETSE_AHBooOlI
&
~
CORETSE_AHBloOlI
}
}
&
CORETSE_AHBOiOlI
[
9
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOiOlI
<=
#
CORETSE_AHBIoII
10
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOiOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBioOlI
[
9
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIiOlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIiOlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOi
;
end
assign
CORETSE_AHBliOlI
=
(
CORETSE_AHBiilOI
&
CORETSE_AHBiiiII
[
3
:
0
]
==
4
'h
3
|
CORETSE_AHBiilOI
&
CORETSE_AHBiiiII
[
3
:
0
]
==
4
'h
1
|
CORETSE_AHBolo
&
CORETSE_AHBoo01
[
1
]
&
~
CORETSE_AHBOIi
&
~
CORETSE_AHBO0o
|
CORETSE_AHBiloII
&
~
CORETSE_AHBoo01
[
1
]
&
~
CORETSE_AHBOIi
&
~
CORETSE_AHBO0o
)
&
~
CORETSE_AHBilo
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBolo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBolo
<=
#
CORETSE_AHBIoII
CORETSE_AHBliOlI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIOIlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIOIlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBolo
;
end
assign
CORETSE_AHBoiOlI
=
CORETSE_AHBiloII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBO0oII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBI1oII
&
~
CORETSE_AHBOliII
&
CORETSE_AHBlIiII
|
CORETSE_AHBOOo1
&
~
CORETSE_AHBiOi
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOOo1
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiOlI
;
end
assign
CORETSE_AHBO0llI
=
CORETSE_AHBiloII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBO0oII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBI1oII
&
~
CORETSE_AHBOliII
&
CORETSE_AHBlIiII
|
CORETSE_AHBI0llI
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBI0llI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBI0llI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0llI
;
end
assign
CORETSE_AHBiiOlI
=
~
CORETSE_AHBO0o
&
CORETSE_AHBoIiII
&
~
CORETSE_AHBii0OI
&
~
CORETSE_AHBOiIlI
&
CORETSE_AHBllOlI
&
~
CORETSE_AHBl0OlI
|
CORETSE_AHBO0o
&
~
(
CORETSE_AHBiOi
&
~
CORETSE_AHBIiOlI
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBO0o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiOlI
;
end
assign
CORETSE_AHBOOIlI
=
CORETSE_AHBOiIlI
|
CORETSE_AHBoIiII
&
CORETSE_AHBllOlI
&
CORETSE_AHBl0OlI
|
CORETSE_AHBoIiII
&
~
CORETSE_AHBllOlI
|
CORETSE_AHBii0OI
|
CORETSE_AHBoIllI
|
CORETSE_AHBilo
&
~
CORETSE_AHBiOi
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBilo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBilo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOIlI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBI0o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBI0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIlOlI
;
end
assign
CORETSE_AHBillII
=
CORETSE_AHBiilOI
|
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
|
CORETSE_AHBl0oII
|
CORETSE_AHBI1oII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBO0lII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBO0lII
<=
#
CORETSE_AHBIoII
CORETSE_AHBillII
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBI0Io
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBI0Io
<=
#
CORETSE_AHBIoII
CORETSE_AHBillII
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBiIIlI
<=
#
CORETSE_AHBIoII
8
'b
0
;
CORETSE_AHBOlIlI
<=
#
CORETSE_AHBIoII
8
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBiIIlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIIlI
;
CORETSE_AHBOlIlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIlIlI
;
end
end
assign
CORETSE_AHBoOIlI
[
7
:
0
]
=
{
8
{
CORETSE_AHBiilOI
}
}
&
{
{
4
{
CORETSE_AHBoo01
[
1
]
}
}
&
{
CORETSE_AHBOO0OI
,
3
'h
5
}
,
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOO0OI
,
3
'h
5
}
|
{
8
{
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
}
}
&
{
CORETSE_AHBiio
[
7
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiOIlI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiOIlI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOIlI
[
7
:
0
]
;
end
generate
if
(
CORETSE_AHBiOI
==
1
)
begin
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlollI
[
9
:
0
]
<=
10
'b
0000000001
;
else
if
(
CORETSE_AHBo1Oo
&
CORETSE_AHBOoo1
&
(
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBOo1II
)
)
CORETSE_AHBlollI
[
9
:
0
]
<=
{
CORETSE_AHBlollI
[
8
:
0
]
,
CORETSE_AHBlollI
[
9
]
}
;
else
CORETSE_AHBlollI
[
9
:
0
]
<=
CORETSE_AHBlollI
[
9
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOo1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOo1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBOio1
;
end
assign
CORETSE_AHBIo1II
=
CORETSE_AHBIoo1
&
CORETSE_AHBOio1
;
assign
CORETSE_AHBIIIlI
=
{
8
{
CORETSE_AHBooo1
}
}
&
CORETSE_AHBiOIlI
|
{
8
{
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
}
}
&
CORETSE_AHBloo1
[
7
:
0
]
|
{
8
{
~
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
}
}
&
CORETSE_AHBiOIlI
;
assign
CORETSE_AHBoIIlI
=
{
8
{
CORETSE_AHBooo1
}
}
&
CORETSE_AHBlIIlI
|
{
8
{
CORETSE_AHBlollI
[
9
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
7
:
0
]
|
{
8
{
CORETSE_AHBlollI
[
8
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
15
:
8
]
|
{
8
{
CORETSE_AHBlollI
[
7
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
23
:
16
]
|
{
8
{
CORETSE_AHBlollI
[
6
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
31
:
24
]
|
{
8
{
CORETSE_AHBlollI
[
5
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
39
:
32
]
|
{
8
{
CORETSE_AHBlollI
[
4
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
47
:
40
]
|
{
8
{
CORETSE_AHBlollI
[
3
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
55
:
48
]
|
{
8
{
CORETSE_AHBlollI
[
2
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
63
:
56
]
|
{
8
{
CORETSE_AHBlollI
[
1
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
71
:
64
]
|
{
8
{
CORETSE_AHBlollI
[
0
]
&
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBioo1
[
79
:
72
]
|
{
8
{
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBloo1
[
15
:
8
]
|
{
8
{
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
~
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBloo1
[
7
:
0
]
|
{
8
{
~
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
~
CORETSE_AHBOoo1
}
}
&
CORETSE_AHBlIIlI
;
assign
CORETSE_AHBIlIlI
=
{
8
{
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
~
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBloo1
[
15
:
8
]
|
{
8
{
~
(
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
~
CORETSE_AHBoo01
[
1
]
)
}
}
&
CORETSE_AHBiIIlI
;
assign
CORETSE_AHBllIlI
=
{
8
{
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
~
CORETSE_AHBoo01
[
1
]
}
}
&
CORETSE_AHBloo1
[
15
:
8
]
|
{
8
{
~
(
CORETSE_AHBIo1II
&
~
CORETSE_AHBooo1
&
~
CORETSE_AHBoo01
[
1
]
)
}
}
&
CORETSE_AHBOlIlI
;
end
else
begin
assign
CORETSE_AHBIIIlI
=
CORETSE_AHBiOIlI
;
assign
CORETSE_AHBoIIlI
=
CORETSE_AHBlIIlI
;
assign
CORETSE_AHBIlIlI
=
CORETSE_AHBiIIlI
;
assign
CORETSE_AHBllIlI
=
CORETSE_AHBOlIlI
;
always
@
(
*
)
CORETSE_AHBlollI
=
10
'b
0
;
end
endgenerate
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlIIlI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBlIIlI
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIIlI
[
7
:
0
]
;
end
assign
CORETSE_AHBI11OI
=
CORETSE_AHBiilOI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBil1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBolIlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBilIlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBil1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBI11OI
;
CORETSE_AHBolIlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBil1o
;
CORETSE_AHBilIlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0IlI
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBlioII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBlioII
<=
#
CORETSE_AHBIoII
CORETSE_AHBolIlI
;
end
end
assign
CORETSE_AHBi0IlI
=
CORETSE_AHBlioII
;
assign
CORETSE_AHBl11OI
=
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
&
CORETSE_AHBoo01
[
1
]
|
CORETSE_AHBl0oII
&
(
CORETSE_AHBoo01
[
1
]
|
~
CORETSE_AHBi0oII
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBol1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBO0IlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBI0IlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBol1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBl11OI
;
CORETSE_AHBO0IlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol1o
;
CORETSE_AHBI0IlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1IlI
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBoioII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBoioII
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0IlI
;
end
end
assign
CORETSE_AHBO1IlI
=
CORETSE_AHBoioII
;
assign
CORETSE_AHBo11OI
=
~
CORETSE_AHBI11OI
&
~
CORETSE_AHBl11OI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBO01o
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBl0IlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBo0IlI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBO01o
<=
#
CORETSE_AHBIoII
CORETSE_AHBo11OI
;
CORETSE_AHBl0IlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO01o
;
CORETSE_AHBo0IlI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1IlI
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBiioII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBiioII
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0IlI
;
end
end
assign
CORETSE_AHBI1IlI
=
CORETSE_AHBiioII
;
pecrc
CORETSE_AHBi1oOI
(
.CORETSE_AHBOl1o
(
CORETSE_AHBiOO1
)
,
.CORETSE_AHBIl1o
(
CORETSE_AHBIio1
)
,
.CORETSE_AHBll1o
(
CORETSE_AHBllIlI
)
,
.CORETSE_AHBol1o
(
CORETSE_AHBI0IlI
)
,
.CORETSE_AHBil1o
(
CORETSE_AHBilIlI
)
,
.CORETSE_AHBO01o
(
CORETSE_AHBo0IlI
)
,
.CORETSE_AHBI01o
(
CORETSE_AHBo1Oo
)
,
.CORETSE_AHBl01o
(
CORETSE_AHBl01o
)
,
.CORETSE_AHBo01o
(
CORETSE_AHBo01o
)
)
;
assign
CORETSE_AHBl1IlI
[
7
:
0
]
=
{
~
CORETSE_AHBl01o
[
24
]
,
~
CORETSE_AHBl01o
[
25
]
,
~
CORETSE_AHBl01o
[
26
]
,
~
CORETSE_AHBl01o
[
27
]
,
~
CORETSE_AHBl01o
[
28
]
,
~
CORETSE_AHBl01o
[
29
]
,
~
CORETSE_AHBl01o
[
30
]
,
~
CORETSE_AHBl01o
[
31
]
}
;
assign
CORETSE_AHBo1IlI
[
7
:
0
]
=
{
~
CORETSE_AHBl01o
[
16
]
,
~
CORETSE_AHBl01o
[
17
]
,
~
CORETSE_AHBl01o
[
18
]
,
~
CORETSE_AHBl01o
[
19
]
,
~
CORETSE_AHBl01o
[
20
]
,
~
CORETSE_AHBl01o
[
21
]
,
~
CORETSE_AHBl01o
[
22
]
,
~
CORETSE_AHBl01o
[
23
]
}
;
assign
CORETSE_AHBi1IlI
[
7
:
0
]
=
{
~
CORETSE_AHBl01o
[
8
]
,
~
CORETSE_AHBl01o
[
9
]
,
~
CORETSE_AHBl01o
[
10
]
,
~
CORETSE_AHBl01o
[
11
]
,
~
CORETSE_AHBl01o
[
12
]
,
~
CORETSE_AHBl01o
[
13
]
,
~
CORETSE_AHBl01o
[
14
]
,
~
CORETSE_AHBl01o
[
15
]
}
;
assign
CORETSE_AHBOoIlI
[
7
:
0
]
=
{
~
CORETSE_AHBl01o
[
0
]
,
~
CORETSE_AHBl01o
[
1
]
,
~
CORETSE_AHBl01o
[
2
]
,
~
CORETSE_AHBl01o
[
3
]
,
~
CORETSE_AHBl01o
[
4
]
,
~
CORETSE_AHBl01o
[
5
]
,
~
CORETSE_AHBl01o
[
6
]
,
~
CORETSE_AHBl01o
[
7
]
}
;
assign
CORETSE_AHBIoIlI
=
CORETSE_AHBO0lII
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBi01II
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBO11II
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBoI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBi01II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoIlI
;
CORETSE_AHBO11II
<=
#
CORETSE_AHBIoII
CORETSE_AHBI11II
;
CORETSE_AHBoI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo1II
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBIOiII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBIOiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBi01II
;
end
end
assign
CORETSE_AHBI11II
=
CORETSE_AHBIOiII
;
assign
CORETSE_AHBloIlI
[
7
:
0
]
=
{
8
{
CORETSE_AHBoo01
[
1
]
&
~|
CORETSE_AHBOIiII
}
}
&
CORETSE_AHBllIlI
[
7
:
0
]
|
{
8
{
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
3
]
}
}
&
(
CORETSE_AHBl1IlI
[
7
:
0
]
^
CORETSE_AHBoliII
)
|
{
8
{
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
2
]
}
}
&
(
CORETSE_AHBo1IlI
[
7
:
0
]
^
CORETSE_AHBoliII
)
|
{
8
{
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
1
]
}
}
&
(
CORETSE_AHBi1IlI
[
7
:
0
]
^
CORETSE_AHBoliII
)
|
{
8
{
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
0
]
}
}
&
(
CORETSE_AHBOoIlI
[
7
:
0
]
^
CORETSE_AHBoliII
)
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
~|
CORETSE_AHBOIiII
&
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
CORETSE_AHBllIlI
[
3
:
0
]
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
~|
CORETSE_AHBOIiII
&
~
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
CORETSE_AHBllIlI
[
7
:
4
]
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
3
]
&
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBl1IlI
[
3
:
0
]
^
CORETSE_AHBoliII
[
3
:
0
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
3
]
&
~
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBl1IlI
[
7
:
4
]
^
CORETSE_AHBoliII
[
7
:
4
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
2
]
&
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBo1IlI
[
3
:
0
]
^
CORETSE_AHBoliII
[
3
:
0
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
2
]
&
~
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBo1IlI
[
7
:
4
]
^
CORETSE_AHBoliII
[
7
:
4
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
1
]
&
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBi1IlI
[
3
:
0
]
^
CORETSE_AHBoliII
[
3
:
0
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
1
]
&
~
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBi1IlI
[
7
:
4
]
^
CORETSE_AHBoliII
[
7
:
4
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
0
]
&
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBOoIlI
[
3
:
0
]
^
CORETSE_AHBoliII
[
3
:
0
]
)
}
|
{
8
{
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBOIiII
[
0
]
&
~
CORETSE_AHBlooII
}
}
&
{
4
'h
0
,
(
CORETSE_AHBOoIlI
[
7
:
4
]
^
CORETSE_AHBoliII
[
7
:
4
]
)
}
;
assign
CORETSE_AHBooIlI
=
CORETSE_AHBloIlI
;
assign
CORETSE_AHBoo1II
=
CORETSE_AHBo11II
;
assign
CORETSE_AHBlo1II
=
CORETSE_AHBO11II
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBII
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBII
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBooIlI
[
7
:
0
]
;
end
assign
CORETSE_AHBioIlI
=
CORETSE_AHBIOllI
|
CORETSE_AHBOOllI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBl11II
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBo11II
<=
#
CORETSE_AHBIoII
1
'b
0
;
CORETSE_AHBOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBl11II
<=
#
CORETSE_AHBIoII
CORETSE_AHBioIlI
;
CORETSE_AHBo11II
<=
#
CORETSE_AHBIoII
CORETSE_AHBi11II
;
CORETSE_AHBOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo1II
;
end
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
begin
CORETSE_AHBOOiII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
else
if
(
CORETSE_AHBo1Oo
)
begin
CORETSE_AHBOOiII
<=
#
CORETSE_AHBIoII
CORETSE_AHBl11II
;
end
end
assign
CORETSE_AHBi11II
=
CORETSE_AHBOOiII
;
assign
CORETSE_AHBIiIlI
=
~
CORETSE_AHBlOllI
&
CORETSE_AHBOliII
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
&
CORETSE_AHBllOlI
&
CORETSE_AHBl0OlI
|
CORETSE_AHBlOllI
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlOllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBlOllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIiIlI
;
end
assign
CORETSE_AHBliIlI
=
~
CORETSE_AHBoOllI
&
CORETSE_AHBoIiII
&
CORETSE_AHBlOoII
&
~
CORETSE_AHBllOlI
|
CORETSE_AHBoOllI
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBoOllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoOllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBliIlI
;
end
assign
CORETSE_AHBii0OI
=
(
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
|
CORETSE_AHBI1oII
)
&
~
CORETSE_AHBIIi
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBIIOlI
;
assign
CORETSE_AHBoiIlI
=
~
CORETSE_AHBOOllI
&
CORETSE_AHBii0OI
|
CORETSE_AHBOOllI
&
~
CORETSE_AHBo1llI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOOllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOOllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiIlI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiOllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiOllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOllI
;
end
assign
CORETSE_AHBOiIlI
=
(
CORETSE_AHBiloII
|
CORETSE_AHBO0oII
)
&
CORETSE_AHBIIi
&
~
CORETSE_AHBlOoII
;
assign
CORETSE_AHBiiIlI
=
~
CORETSE_AHBIOllI
&
CORETSE_AHBOiIlI
|
CORETSE_AHBIOllI
&
~
CORETSE_AHBo1llI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIOllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIOllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiIlI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOIllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOIllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOllI
;
end
assign
CORETSE_AHBIIllI
=
~
CORETSE_AHBoOi1
&
CORETSE_AHBiIoII
&
CORETSE_AHBiOi
&
(
CORETSE_AHBoo01
[
1
:
0
]
==
2
'b
01
&
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
17b7
|
CORETSE_AHBoo01
[
1
:
0
]
==
2
'b
10
&
CORETSE_AHBoOOlI
[
15
:
0
]
==
16
'h
0bdb
)
|
CORETSE_AHBoOi1
&
~
CORETSE_AHBIOo1
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBoOi1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoOi1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIllI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOlllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOlllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIllI
&
~
CORETSE_AHBoOi1
;
end
assign
CORETSE_AHBlIllI
=
~
CORETSE_AHBoIllI
&
CORETSE_AHBOlllI
&
~
CORETSE_AHBloi1
|
CORETSE_AHBoIllI
&
~
CORETSE_AHBo1llI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBoIllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBoIllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIllI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiIllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiIllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIllI
;
end
assign
CORETSE_AHBolllI
=
~
CORETSE_AHBlOllI
&
~
CORETSE_AHBoOllI
&
~
CORETSE_AHBOOllI
&
~
CORETSE_AHBIOllI
&
~
CORETSE_AHBoIllI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBilllI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBilllI
<=
#
CORETSE_AHBIoII
CORETSE_AHBolllI
;
end
assign
CORETSE_AHBIo1OI
=
CORETSE_AHBil0OI
&
CORETSE_AHBIOIlI
&
CORETSE_AHBOIIlI
[
0
]
|
~
(
CORETSE_AHBil0OI
&
CORETSE_AHBIOIlI
)
&
CORETSE_AHBOl00
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOl00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOl00
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo1OI
;
end
assign
CORETSE_AHBlo1OI
=
CORETSE_AHBil0OI
&
CORETSE_AHBIOIlI
&
(
&
CORETSE_AHBOIIlI
[
7
:
0
]
)
|
CORETSE_AHBO00OI
&
CORETSE_AHBIOIlI
&
(
&
CORETSE_AHBOIIlI
[
7
:
0
]
)
&
CORETSE_AHBiI00
|
CORETSE_AHBI00OI
&
CORETSE_AHBIOIlI
&
(
&
CORETSE_AHBOIIlI
[
7
:
0
]
)
&
CORETSE_AHBiI00
|
CORETSE_AHBl00OI
&
CORETSE_AHBIOIlI
&
(
&
CORETSE_AHBOIIlI
[
7
:
0
]
)
&
CORETSE_AHBiI00
|
CORETSE_AHBo00OI
&
CORETSE_AHBIOIlI
&
(
&
CORETSE_AHBOIIlI
[
7
:
0
]
)
&
CORETSE_AHBiI00
|
CORETSE_AHBO10OI
&
CORETSE_AHBIOIlI
&
(
&
CORETSE_AHBOIIlI
[
7
:
0
]
)
&
CORETSE_AHBiI00
|
(
CORETSE_AHBOIOlI
|
~
CORETSE_AHBIOIlI
)
&
CORETSE_AHBiI00
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBiI00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBiI00
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo1OI
;
end
assign
CORETSE_AHBoo1OI
=
CORETSE_AHBl10OI
&
CORETSE_AHBIOIlI
|
CORETSE_AHBOo0OI
&
CORETSE_AHBIOIlI
&
CORETSE_AHBOOoOI
;
assign
CORETSE_AHBio1OI
=
CORETSE_AHBo1oOI
&
CORETSE_AHBIOIlI
|
CORETSE_AHBiOOlI
&
CORETSE_AHBIOIlI
&
CORETSE_AHBOOoOI
;
assign
CORETSE_AHBOi1OI
[
15
:
0
]
=
{
16
{
CORETSE_AHBoo1OI
}
}
&
{
CORETSE_AHBOIIlI
[
7
:
0
]
,
CORETSE_AHBIi1OI
[
7
:
0
]
}
|
{
16
{
CORETSE_AHBio1OI
}
}
&
{
CORETSE_AHBIi1OI
[
15
:
8
]
,
CORETSE_AHBOIIlI
[
7
:
0
]
}
|
{
16
{
~
CORETSE_AHBoo1OI
&
~
CORETSE_AHBio1OI
}
}
&
{
CORETSE_AHBIi1OI
[
15
:
8
]
,
CORETSE_AHBIi1OI
[
7
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIi1OI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBIi1OI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi1OI
[
15
:
0
]
;
end
assign
CORETSE_AHBli1OI
=
CORETSE_AHBIi1OI
[
15
:
0
]
>
16
'h
05dc
;
assign
CORETSE_AHBoi1OI
=
(
CORETSE_AHBIi1OI
[
15
:
0
]
>=
16
'h
002e
&
~
CORETSE_AHBOOoOI
|
CORETSE_AHBIi1OI
[
15
:
0
]
>=
16
'h
002a
&
CORETSE_AHBOOoOI
)
;
assign
CORETSE_AHBl0llI
=
(
CORETSE_AHBiOoOI
[
15
:
0
]
>=
16
'h
002e
&
~
CORETSE_AHBOOoOI
|
CORETSE_AHBiOoOI
[
15
:
0
]
>=
16
'h
002a
&
CORETSE_AHBOOoOI
)
;
assign
CORETSE_AHBii1OI
=
CORETSE_AHBo10OI
&
CORETSE_AHBIOIlI
&
CORETSE_AHBIi1OI
[
15
:
0
]
==
16
'h
8100
|
(
~
CORETSE_AHBo10OI
|
~
CORETSE_AHBIOIlI
)
&
CORETSE_AHBOOoOI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOOoOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBOOoOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1OI
;
end
assign
CORETSE_AHBo0llI
=
CORETSE_AHBli1OI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBi0llI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi0llI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0llI
;
end
assign
CORETSE_AHBiOoOI
=
{
16
{
~
CORETSE_AHBOOoOI
}
}
&
(
CORETSE_AHBoOOlI
[
15
:
0
]
-
5
'h
12
)
|
{
16
{
CORETSE_AHBOOoOI
}
}
&
(
CORETSE_AHBoOOlI
[
15
:
0
]
-
5
'h
16
)
;
assign
CORETSE_AHBO1llI
=
CORETSE_AHBoo01
[
0
]
&
(
CORETSE_AHBIi1OI
[
15
:
0
]
!=
CORETSE_AHBiOoOI
[
15
:
0
]
+
1
)
|
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBIi1OI
[
15
:
0
]
!=
CORETSE_AHBiOoOI
[
15
:
0
]
;
assign
CORETSE_AHBOIoOI
=
CORETSE_AHBi0i1
&
(
CORETSE_AHBoi1OI
&
~
CORETSE_AHBli1OI
&
CORETSE_AHBO1llI
|
~
CORETSE_AHBoi1OI
&
CORETSE_AHBl0llI
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIIoOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIIoOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIoOI
;
end
assign
CORETSE_AHBI1llI
=
~
CORETSE_AHBo1llI
&
(
CORETSE_AHBiloII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBO0oII
&
~
CORETSE_AHBlOoII
&
CORETSE_AHBOIi
&
~
(
CORETSE_AHBlIoII
|
CORETSE_AHBIIoII
)
|
CORETSE_AHBI1oII
&
~
CORETSE_AHBOliII
&
CORETSE_AHBlIiII
|
CORETSE_AHBOliII
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
&
CORETSE_AHBllOlI
&
CORETSE_AHBl0OlI
|
CORETSE_AHBoOllI
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
&
~
CORETSE_AHBllOlI
|
CORETSE_AHBOOllI
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
|
CORETSE_AHBIOllI
&
CORETSE_AHBI1oII
&
CORETSE_AHBlIiII
|
CORETSE_AHBoIllI
&
CORETSE_AHBiIllI
&
CORETSE_AHBlIllI
)
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBo1llI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBo1llI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1llI
;
end
assign
CORETSE_AHBl1llI
=
CORETSE_AHBo1llI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBi1llI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBi1llI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1llI
;
end
assign
CORETSE_AHBOollI
=
CORETSE_AHBi1llI
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBIOo1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBIOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOollI
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBOi1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
&
CORETSE_AHBiOi
&
CORETSE_AHBolo
)
CORETSE_AHBOi1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBilIo
;
else
if
(
CORETSE_AHBo1Oo
&
CORETSE_AHBIOo1
)
CORETSE_AHBOi1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOi1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi1II
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBio1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBo1Oo
&
CORETSE_AHBiOi
&
CORETSE_AHBolo
)
CORETSE_AHBio1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOo1
;
else
if
(
CORETSE_AHBo1Oo
&
CORETSE_AHBIOo1
)
CORETSE_AHBio1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBio1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBio1II
;
end
assign
CORETSE_AHBIollI
[
51
:
48
]
=
{
4
{
CORETSE_AHBi1llI
}
}
&
{
CORETSE_AHBOOoOI
,
CORETSE_AHBllllI
,
CORETSE_AHBOi1II
,
CORETSE_AHBio1II
}
|
{
4
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
51
:
48
]
;
assign
CORETSE_AHBIollI
[
47
:
32
]
=
{
16
{
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBOlOlI
[
15
:
0
]
|
{
16
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
47
:
32
]
;
assign
CORETSE_AHBIollI
[
31
:
28
]
=
{
4
{
CORETSE_AHBi1llI
}
}
&
{
CORETSE_AHBOIllI
,
CORETSE_AHBiOllI
,
CORETSE_AHBoOllI
,
CORETSE_AHBlOllI
}
|
{
4
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
31
:
28
]
;
assign
CORETSE_AHBIollI
[
27
:
24
]
=
{
4
{
CORETSE_AHBi1llI
}
}
&
{
CORETSE_AHBoOi1
,
CORETSE_AHBilllI
&
CORETSE_AHBi0iII
,
CORETSE_AHBilllI
&
CORETSE_AHBiI00
,
CORETSE_AHBilllI
&
CORETSE_AHBOl00
}
|
{
4
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
27
:
24
]
;
assign
CORETSE_AHBIollI
[
23
:
20
]
=
{
4
{
CORETSE_AHBi1llI
}
}
&
{
CORETSE_AHBilllI
&
CORETSE_AHBI0llI
,
CORETSE_AHBilllI
&
CORETSE_AHBi0llI
,
CORETSE_AHBilllI
&
CORETSE_AHBIIoOI
,
CORETSE_AHBilllI
&
~
CORETSE_AHBo1oII
&
CORETSE_AHBo01o
}
|
{
4
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
23
:
20
]
;
assign
CORETSE_AHBIollI
[
19
:
16
]
=
{
4
{
CORETSE_AHBi1llI
}
}
&
{
4
{
CORETSE_AHBilllI
}
}
&
CORETSE_AHBI0OlI
[
3
:
0
]
|
{
4
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
19
:
16
]
;
assign
CORETSE_AHBIollI
[
15
:
0
]
=
{
16
{
CORETSE_AHBi1llI
}
}
&
{
16
{
CORETSE_AHBilllI
}
}
&
CORETSE_AHBoOOlI
[
15
:
0
]
|
{
16
{
~
CORETSE_AHBi1llI
}
}
&
CORETSE_AHBlOo1
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBIio1
)
begin
if
(
CORETSE_AHBIio1
)
CORETSE_AHBlOo1
<=
#
CORETSE_AHBIoII
52
'h
0
;
else
if
(
CORETSE_AHBo1Oo
)
CORETSE_AHBlOo1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIollI
[
51
:
0
]
;
end
endmodule
