module
CoreTSE_Webserver_CORETSE_AHB_0_CORETSE_AHB
(
STBP
,
TXCLK
,
RXCLK
,
GTXCLK
,
PMARX_CLK0
,
PMARX_CLK1
,
RCG
,
TCG
,
SIGNAL_DETECT
,
TXD
,
TXEN
,
TXER
,
RXD
,
RXDV
,
RXER
,
CRS
,
COL
,
HRESETN
,
HCLK
,
HREADY
,
HWDATA
,
HADDR
,
HSEL
,
HTRANS
,
HWRITE
,
HRDATA
,
HRESP
,
HREADYOUT
,
HBURST
,
HMASTLOCK
,
HSIZE
,
TXHGRANT
,
TXHRESP
,
TXHRDATA
,
TXHBUSREQ
,
TXHTRANS
,
TXHADDR
,
TXHWRITE
,
TXHWDATA
,
TXHREADY
,
TXHBURST
,
TXHLOCK
,
TXHSIZE
,
RXHGRANT
,
RXHRESP
,
RXHRDATA
,
RXHBUSREQ
,
RXHTRANS
,
RXHADDR
,
RXHWRITE
,
RXHWDATA
,
RXHREADY
,
RXHBURST
,
RXHLOCK
,
RXHSIZE
,
MDI
,
MDC
,
MDO
,
MDOEN
,
TBI_READY
,
TBI_TXVAL
,
TSM_CONTROL
,
TSM_INTR
,
ANX_STATE
,
SYNC
)
;
parameter
FAMILY
=
19
;
parameter
GMII_TBI
=
0
;
parameter
PACKET_SIZE
=
11
;
parameter
SAL
=
1
;
parameter
WOL
=
1
;
parameter
STATS
=
1
;
parameter
MDIO_PHYID
=
18
;
input
STBP
;
input
TXCLK
;
input
RXCLK
;
input
GTXCLK
;
input
PMARX_CLK0
;
input
PMARX_CLK1
;
input
[
9
:
0
]
RCG
;
output
[
9
:
0
]
TCG
;
input
SIGNAL_DETECT
;
output
[
7
:
0
]
TXD
;
output
TXEN
;
output
TXER
;
input
[
7
:
0
]
RXD
;
input
RXDV
;
input
RXER
;
input
CRS
;
input
COL
;
input
HRESETN
;
input
HCLK
;
input
HSEL
;
input
[
31
:
0
]
HADDR
;
input
HWRITE
;
input
[
1
:
0
]
HTRANS
;
input
[
2
:
0
]
HSIZE
;
input
[
2
:
0
]
HBURST
;
input
HMASTLOCK
;
input
HREADY
;
input
[
31
:
0
]
HWDATA
;
output
HREADYOUT
;
output
[
1
:
0
]
HRESP
;
output
[
31
:
0
]
HRDATA
;
input
TXHGRANT
;
input
TXHREADY
;
input
[
1
:
0
]
TXHRESP
;
input
[
31
:
0
]
TXHRDATA
;
output
TXHBUSREQ
;
output
TXHLOCK
;
output
[
1
:
0
]
TXHTRANS
;
output
[
31
:
0
]
TXHADDR
;
output
TXHWRITE
;
output
[
2
:
0
]
TXHSIZE
;
output
[
2
:
0
]
TXHBURST
;
output
[
31
:
0
]
TXHWDATA
;
input
RXHGRANT
;
input
RXHREADY
;
input
[
1
:
0
]
RXHRESP
;
input
[
31
:
0
]
RXHRDATA
;
output
RXHBUSREQ
;
output
RXHLOCK
;
output
[
1
:
0
]
RXHTRANS
;
output
[
31
:
0
]
RXHADDR
;
output
RXHWRITE
;
output
[
2
:
0
]
RXHSIZE
;
output
[
2
:
0
]
RXHBURST
;
output
[
31
:
0
]
RXHWDATA
;
input
MDI
;
output
MDC
;
output
MDO
;
output
MDOEN
;
output
[
31
:
0
]
TSM_CONTROL
;
output
[
2
:
0
]
TSM_INTR
;
input
TBI_READY
;
output
TBI_TXVAL
;
output
[
9
:
0
]
ANX_STATE
;
output
SYNC
;
CoreTSE_top
#
(
.FAMILY
(
FAMILY
)
,
.GMII_TBI
(
GMII_TBI
)
,
.MCXMAC_SAL_ON
(
SAL
)
,
.MCXMAC_STATS_ON
(
STATS
)
,
.MCXMAC_WOL_ON
(
WOL
)
,
.MDIO_PHYID
(
MDIO_PHYID
)
,
.RABITS
(
(
PACKET_SIZE
+
1
)
)
,
.TABITS
(
PACKET_SIZE
)
)
CoreTSE_top_inst
(
.RSTBP_I
(
STBP
)
,
.TXCLK_I
(
TXCLK
)
,
.RXCLK_I
(
RXCLK
)
,
.GTXCLK_I
(
GTXCLK
)
,
.PMARX_CLK0_I
(
PMARX_CLK0
)
,
.PMARX_CLK1_I
(
PMARX_CLK1
)
,
.TSMAC_RCG_I
(
RCG
)
,
.TSMAC_RXD_I
(
RXD
)
,
.TSMAC_RXDV_I
(
RXDV
)
,
.TSMAC_RXER_I
(
RXER
)
,
.TSMAC_CRS_I
(
CRS
)
,
.TSMAC_COL_I
(
COL
)
,
.HRESET_NI
(
HRESETN
)
,
.HCLK_I
(
HCLK
)
,
.AHBS_HREADY_I
(
HREADY
)
,
.AHBS_HWDATA_I
(
HWDATA
)
,
.AHBS_HADDR_I
(
HADDR
)
,
.AHBS_HSEL_I
(
HSEL
)
,
.AHBS_HTRANS_I
(
HTRANS
)
,
.AHBS_HWRITE_I
(
HWRITE
)
,
.AHBS_HBURST_I
(
HBURST
[
0
]
)
,
.AHBS_HMASTLOCK_I
(
HMASTLOCK
)
,
.AHBS_HPROT_I
(
)
,
.AHBS_HSIZE_I
(
HSIZE
[
0
]
)
,
.AHBM_TXHGRANT_I
(
TXHGRANT
)
,
.AHBM_TXHRESPM_I
(
TXHRESP
)
,
.AHBM_TXHRDATAM_I
(
TXHRDATA
)
,
.AHBM_TXHREADY_I
(
TXHREADY
)
,
.AHBM_RXHGRANT_I
(
RXHGRANT
)
,
.AHBM_RXHRESPM_I
(
RXHRESP
)
,
.AHBM_RXHRDATAM_I
(
RXHRDATA
)
,
.AHBM_RXHREADY_I
(
RXHREADY
)
,
.MGMT_MDI_I
(
MDI
)
,
.TBI_READY_I
(
TBI_READY
)
,
.SIGNAL_DETECT_I
(
SIGNAL_DETECT
)
,
.TSMAC_TCG_O
(
TCG
)
,
.TSMAC_TXD_O
(
TXD
)
,
.TSMAC_TXEN_O
(
TXEN
)
,
.TSMAC_TXER_O
(
TXER
)
,
.AHBS_HRDATA_O
(
HRDATA
)
,
.AHBS_HRESP_O
(
HRESP
)
,
.AHBS_HREADY_O
(
HREADYOUT
)
,
.AHBM_TXHBUSREQ_O
(
TXHBUSREQ
)
,
.AHBM_TXHTRANSM_O
(
TXHTRANS
)
,
.AHBM_TXHADDRM_O
(
TXHADDR
)
,
.AHBM_TXHWRITEM_O
(
TXHWRITE
)
,
.AHBM_TXHWDATAM_O
(
TXHWDATA
)
,
.AHBM_RXHBUSREQ_O
(
RXHBUSREQ
)
,
.AHBM_RXHTRANSM_O
(
RXHTRANS
)
,
.AHBM_RXHADDRM_O
(
RXHADDR
)
,
.AHBM_RXHWRITEM_O
(
RXHWRITE
)
,
.AHBM_RXHWDATAM_O
(
RXHWDATA
)
,
.AHBM_TXHBURST_O
(
TXHBURST
)
,
.AHBM_RXHBURST_O
(
RXHBURST
)
,
.AHBM_TXMASTLOCK_O
(
CORETSE_AHBO
)
,
.AHBM_RXMASTLOCK_O
(
CORETSE_AHBI
)
,
.AHBM_TXHSIZE_O
(
TXHSIZE
)
,
.AHBM_RXHSIZE_O
(
RXHSIZE
)
,
.AHBM_TXHSPLIT_O
(
)
,
.AHBM_RXHSPLIT_O
(
)
,
.AHBM_TXHSEL_O
(
)
,
.AHBM_RXHSEL_O
(
)
,
.MGMT_MDC_O
(
MDC
)
,
.MGMT_MDO_O
(
MDO
)
,
.MGMT_MDOEN_O
(
MDOEN
)
,
.TBI_TXVAL_O
(
TBI_TXVAL
)
,
.TSM_CONTROL_O
(
TSM_CONTROL
)
,
.TSM_INTR_O
(
TSM_INTR
)
,
.ANX_STATE_O
(
ANX_STATE
)
,
.SYNC_O
(
SYNC
)
)
;
endmodule
