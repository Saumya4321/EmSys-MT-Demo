//                        Proprietary and Confidential 
// REVISION    : $Revision: 1.20 $ 
`include "include.v"
module
ptp_top
#
(
parameter
CORETSE_AHBIII
=
1
,
parameter
CORETSE_AHBlII
=
2
,
parameter
CORETSE_AHBoII
=
1
,
parameter
CORETSE_AHBiII
=
2
,
parameter
CORETSE_AHBOlI
=
18
,
parameter
CORETSE_AHBIlI
=
18
,
parameter
CORETSE_AHBllI
=
5
,
parameter
CORETSE_AHBolI
=
5
)
(
input
CORETSE_AHBiil0,
input
CORETSE_AHBi10lI,
input
CORETSE_AHBOl0,
input
CORETSE_AHBOo0lI,
input
CORETSE_AHBl0I,
input
CORETSE_AHBIl0,
input
CORETSE_AHBOI01I,
input
CORETSE_AHBII01I,
input
CORETSE_AHBlI01I,
input
CORETSE_AHBoI01I,
input
[
1
:
0
]
CORETSE_AHBoIo0I,
input
[
7
:
0
]
CORETSE_AHBiI01I,
input
[
7
:
0
]
CORETSE_AHBOl01I,
input
CORETSE_AHBi1O1I,
input
CORETSE_AHBOOo0I,
input
CORETSE_AHBIOo0I,
input
CORETSE_AHBlo0lI,
input
CORETSE_AHBoo0lI,
input
[
4
:
0
]
CORETSE_AHBoO00,
input
[
31
:
0
]
CORETSE_AHBioo1I,
input
CORETSE_AHBiOo0I,
input
[
7
:
0
]
CORETSE_AHBOIo0I,
input
[
7
:
0
]
CORETSE_AHBIIo0I,
input
CORETSE_AHBOoO1I,
input
CORETSE_AHBlIo0I,
input
CORETSE_AHBiIo0I,
input
CORETSE_AHBlI0,
input
CORETSE_AHBoI0,
input
CORETSE_AHBiI0,
output
[
31
:
0
]
CORETSE_AHBOio1I,
output
CORETSE_AHBIio1I,
output
CORETSE_AHBOl1lI,
output
CORETSE_AHBlio1I,
output
CORETSE_AHBO001I,
output
CORETSE_AHBl001I,
output
[
15
:
0
]
CORETSE_AHBo001I,
output
CORETSE_AHBI101I,
output
CORETSE_AHBO101I,
output
[
79
:
0
]
CORETSE_AHBoio1I,
output
CORETSE_AHBll0,
output
CORETSE_AHBol0,
output
CORETSE_AHBil0,
output
CORETSE_AHBO00,
output
CORETSE_AHBI00
)
;
wire
CORETSE_AHBiio1I
;
wire
[
79
:
0
]
CORETSE_AHBiiI1I
;
wire
CORETSE_AHBI1l1I
;
wire
CORETSE_AHBOo01I
;
wire
CORETSE_AHBOOi1I
;
wire
CORETSE_AHBIOi1I
;
wire
CORETSE_AHBlOi1I
;
wire
[
3
:
0
]
CORETSE_AHBoOi1I
;
wire
[
15
:
0
]
CORETSE_AHBiOi1I
;
wire
[
79
:
0
]
CORETSE_AHBOIi1I
;
wire
[
79
:
0
]
CORETSE_AHBIIi1I
;
wire
[
3
:
0
]
CORETSE_AHBlIi1I
;
wire
[
15
:
0
]
CORETSE_AHBoIi1I
;
wire
[
79
:
0
]
CORETSE_AHBiIi1I
;
wire
[
79
:
0
]
CORETSE_AHBOli1I
;
wire
[
79
:
0
]
CORETSE_AHBIli1I
;
wire
[
79
:
0
]
CORETSE_AHBlli1I
;
wire
[
79
:
0
]
CORETSE_AHBoli1I
;
wire
[
7
:
0
]
CORETSE_AHBiiolI
;
wire
[
7
:
0
]
CORETSE_AHBIOilI
;
wire
CORETSE_AHBili1I
;
wire
CORETSE_AHBolI0I
;
wire
CORETSE_AHBoOl1I
;
wire
CORETSE_AHBO0i1I
;
wire
CORETSE_AHBI0i1I
;
wire
CORETSE_AHBl0i1I
;
wire
CORETSE_AHBo0i1I
;
wire
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
CORETSE_AHBi0i1I
;
wire
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
CORETSE_AHBO1i1I
;
wire
CORETSE_AHBI1i1I
;
wire
CORETSE_AHBl1i1I
;
wire
CORETSE_AHBo1i1I
;
wire
CORETSE_AHBi1i1I
;
wire
CORETSE_AHBOoi1I
;
wire
CORETSE_AHBIoi1I
;
wire
CORETSE_AHBloi1I
;
wire
[
`CORETSE_AHBIoI0
:
0
]
CORETSE_AHBIol0I
;
wire
CORETSE_AHBiol1I
;
wire
CORETSE_AHBlll0I
;
assign
CORETSE_AHBoio1I
=
CORETSE_AHBIIi1I
;
ptp_hstinf
#
(
.CORETSE_AHBlII
(
CORETSE_AHBlII
)
,
.CORETSE_AHBIII
(
CORETSE_AHBIII
)
,
.CORETSE_AHBiII
(
CORETSE_AHBiII
)
,
.CORETSE_AHBoII
(
CORETSE_AHBoII
)
,
.CORETSE_AHBOlI
(
CORETSE_AHBOlI
)
,
.CORETSE_AHBIlI
(
CORETSE_AHBIlI
)
,
.CORETSE_AHBllI
(
CORETSE_AHBllI
)
,
.CORETSE_AHBolI
(
CORETSE_AHBolI
)
)
CORETSE_AHBooi1I
(
.CORETSE_AHBiil0
(
CORETSE_AHBiil0
)
,
.CORETSE_AHBi10lI
(
CORETSE_AHBi10lI
)
,
.CORETSE_AHBOl0
(
CORETSE_AHBOl0
)
,
.CORETSE_AHBOo0lI
(
CORETSE_AHBiol1I
)
,
.CORETSE_AHBIo0lI
(
CORETSE_AHBiio1I
)
,
.CORETSE_AHBlo0lI
(
CORETSE_AHBlo0lI
)
,
.CORETSE_AHBoo0lI
(
CORETSE_AHBoo0lI
)
,
.CORETSE_AHBoO00
(
CORETSE_AHBoO00
)
,
.CORETSE_AHBio0lI
(
CORETSE_AHBioo1I
)
,
.CORETSE_AHBOi0lI
(
CORETSE_AHBiiI1I
)
,
.CORETSE_AHBIi0lI
(
CORETSE_AHBI1l1I
)
,
.CORETSE_AHBIl1lI
(
CORETSE_AHBlll0I
)
,
.CORETSE_AHBli0lI
(
CORETSE_AHBOo01I
)
,
.CORETSE_AHBoi0lI
(
CORETSE_AHBOOi1I
)
,
.CORETSE_AHBii0lI
(
CORETSE_AHBIOi1I
)
,
.CORETSE_AHBOO1lI
(
CORETSE_AHBlOi1I
)
,
.CORETSE_AHBIO1lI
(
CORETSE_AHBoOi1I
)
,
.CORETSE_AHBlO1lI
(
CORETSE_AHBiOi1I
)
,
.CORETSE_AHBoO1lI
(
CORETSE_AHBOIi1I
)
,
.CORETSE_AHBioo1
(
CORETSE_AHBIIi1I
)
,
.CORETSE_AHBiO1lI
(
CORETSE_AHBlIi1I
)
,
.CORETSE_AHBOI1lI
(
CORETSE_AHBoIi1I
)
,
.CORETSE_AHBII1lI
(
CORETSE_AHBiIi1I
)
,
.CORETSE_AHBlI1lI
(
CORETSE_AHBOli1I
)
,
.CORETSE_AHBlI0
(
CORETSE_AHBlI0
)
,
.CORETSE_AHBoI0
(
CORETSE_AHBoI0
)
,
.CORETSE_AHBiI0
(
CORETSE_AHBiI0
)
,
.CORETSE_AHBoI1lI
(
CORETSE_AHBOio1I
)
,
.CORETSE_AHBiI1lI
(
CORETSE_AHBIio1I
)
,
.CORETSE_AHBOl1lI
(
CORETSE_AHBOl1lI
)
,
.CORETSE_AHBli1lI
(
CORETSE_AHBlio1I
)
,
.CORETSE_AHBll1lI
(
CORETSE_AHBIli1I
)
,
.CORETSE_AHBol1lI
(
CORETSE_AHBlli1I
)
,
.CORETSE_AHBil1lI
(
CORETSE_AHBoli1I
)
,
.CORETSE_AHBO01lI
(
CORETSE_AHBiiolI
)
,
.CORETSE_AHBI01lI
(
CORETSE_AHBIOilI
)
,
.CORETSE_AHBl01lI
(
CORETSE_AHBili1I
)
,
.CORETSE_AHBo01lI
(
CORETSE_AHBolI0I
)
,
.CORETSE_AHBi01lI
(
CORETSE_AHBoOl1I
)
,
.CORETSE_AHBO11lI
(
CORETSE_AHBO0i1I
)
,
.CORETSE_AHBI11lI
(
CORETSE_AHBI0i1I
)
,
.CORETSE_AHBl11lI
(
CORETSE_AHBl0i1I
)
,
.CORETSE_AHBo11lI
(
CORETSE_AHBo0i1I
)
,
.CORETSE_AHBi11lI
(
CORETSE_AHBloi1I
)
,
.CORETSE_AHBOo1lI
(
CORETSE_AHBIol0I
)
,
.CORETSE_AHBIo1lI
(
CORETSE_AHBi0i1I
)
,
.CORETSE_AHBlo1lI
(
CORETSE_AHBO1i1I
)
,
.CORETSE_AHBoo1lI
(
CORETSE_AHBI1i1I
)
,
.CORETSE_AHBio1lI
(
CORETSE_AHBl1i1I
)
,
.CORETSE_AHBOi1lI
(
CORETSE_AHBo1i1I
)
,
.CORETSE_AHBIi1lI
(
CORETSE_AHBi1i1I
)
,
.CORETSE_AHBoi1lI
(
CORETSE_AHBOoi1I
)
,
.CORETSE_AHBii1lI
(
CORETSE_AHBIoi1I
)
)
;
ptp_tfp
CORETSE_AHBioi1I
(
.CORETSE_AHBOI01I
(
CORETSE_AHBOI01I
)
,
.CORETSE_AHBII01I
(
CORETSE_AHBII01I
)
,
.CORETSE_AHBlOo0I
(
CORETSE_AHBlll0I
)
,
.CORETSE_AHBlI01I
(
CORETSE_AHBlI01I
)
,
.CORETSE_AHBoI01I
(
CORETSE_AHBoI01I
)
,
.CORETSE_AHBoIo0I
(
CORETSE_AHBoIo0I
)
,
.CORETSE_AHBiI01I
(
CORETSE_AHBiI01I
)
,
.CORETSE_AHBOl01I
(
CORETSE_AHBOl01I
)
,
.CORETSE_AHBi1O1I
(
CORETSE_AHBi1O1I
)
,
.CORETSE_AHBIl01I
(
CORETSE_AHBO0i1I
)
,
.CORETSE_AHBoOo0I
(
CORETSE_AHBolI0I
)
,
.CORETSE_AHBll01I
(
CORETSE_AHBIIi1I
)
,
.CORETSE_AHBol01I
(
CORETSE_AHBi1i1I
)
,
.CORETSE_AHBil01I
(
CORETSE_AHBOoi1I
)
,
.CORETSE_AHBO001I
(
CORETSE_AHBO001I
)
,
.CORETSE_AHBIlo0I
(
CORETSE_AHBiOi1I
)
,
.CORETSE_AHBllo0I
(
CORETSE_AHBOIi1I
)
,
.CORETSE_AHBolo0I
(
CORETSE_AHBoOi1I
)
,
.CORETSE_AHBI001I
(
CORETSE_AHBOo01I
)
,
.CORETSE_AHBl001I
(
CORETSE_AHBl001I
)
,
.CORETSE_AHBo001I
(
CORETSE_AHBo001I
)
,
.CORETSE_AHBI101I
(
CORETSE_AHBI101I
)
,
.CORETSE_AHBO101I
(
CORETSE_AHBO101I
)
,
.CORETSE_AHBi001I
(
CORETSE_AHBIOi1I
)
)
;
ptp_rfp
CORETSE_AHBOii1I
(
.CORETSE_AHBOOo0I
(
CORETSE_AHBOOo0I
)
,
.CORETSE_AHBIOo0I
(
CORETSE_AHBIOo0I
)
,
.CORETSE_AHBlOo0I
(
CORETSE_AHBlll0I
)
,
.CORETSE_AHBiOo0I
(
CORETSE_AHBiOo0I
)
,
.CORETSE_AHBoOo0I
(
CORETSE_AHBolI0I
)
,
.CORETSE_AHBOIo0I
(
CORETSE_AHBOIo0I
)
,
.CORETSE_AHBIIo0I
(
CORETSE_AHBIIo0I
)
,
.CORETSE_AHBlIo0I
(
CORETSE_AHBlIo0I
)
,
.CORETSE_AHBiIo0I
(
CORETSE_AHBiIo0I
)
,
.CORETSE_AHBoIo0I
(
CORETSE_AHBoIo0I
)
,
.CORETSE_AHBOlo0I
(
CORETSE_AHBIoi1I
)
,
.CORETSE_AHBIlo0I
(
CORETSE_AHBoIi1I
)
,
.CORETSE_AHBllo0I
(
CORETSE_AHBiIi1I
)
,
.CORETSE_AHBolo0I
(
CORETSE_AHBlIi1I
)
,
.CORETSE_AHBilo0I
(
CORETSE_AHBlOi1I
)
)
;
ptp_rtc
#
(
.CORETSE_AHBlII
(
CORETSE_AHBlII
)
,
.CORETSE_AHBIII
(
CORETSE_AHBIII
)
,
.CORETSE_AHBiII
(
CORETSE_AHBiII
)
,
.CORETSE_AHBoII
(
CORETSE_AHBoII
)
)
CORETSE_AHBIii1I
(
.CORETSE_AHBOl0
(
CORETSE_AHBOl0
)
,
.CORETSE_AHBOo0lI
(
CORETSE_AHBOo0lI
)
,
.CORETSE_AHBl0I
(
CORETSE_AHBl0I
)
,
.CORETSE_AHBlOo0I
(
CORETSE_AHBlll0I
)
,
.CORETSE_AHBIl0
(
CORETSE_AHBIl0
)
,
.CORETSE_AHBilO1I
(
CORETSE_AHBIOilI
)
,
.CORETSE_AHBolO1I
(
CORETSE_AHBiiolI
)
,
.CORETSE_AHBO0O1I
(
CORETSE_AHBl0i1I
)
,
.CORETSE_AHBI0O1I
(
CORETSE_AHBo0i1I
)
,
.CORETSE_AHBl0O1I
(
CORETSE_AHBlli1I
)
,
.CORETSE_AHBo0O1I
(
CORETSE_AHBoli1I
)
,
.CORETSE_AHBloO1I
(
CORETSE_AHBi0i1I
)
,
.CORETSE_AHBooO1I
(
CORETSE_AHBO1i1I
)
,
.CORETSE_AHBoOo0I
(
CORETSE_AHBolI0I
)
,
.CORETSE_AHBi0O1I
(
CORETSE_AHBoOl1I
)
,
.CORETSE_AHBO1O1I
(
CORETSE_AHBloi1I
)
,
.CORETSE_AHBI1O1I
(
CORETSE_AHBIli1I
)
,
.CORETSE_AHBl1O1I
(
CORETSE_AHBili1I
)
,
.CORETSE_AHBo1O1I
(
CORETSE_AHBI0i1I
)
,
.CORETSE_AHBi1O1I
(
CORETSE_AHBi1O1I
)
,
.CORETSE_AHBOoO1I
(
CORETSE_AHBOoO1I
)
,
.CORETSE_AHBIoO1I
(
CORETSE_AHBI1i1I
)
,
.CORETSE_AHBioO1I
(
CORETSE_AHBl1i1I
)
,
.CORETSE_AHBOiO1I
(
CORETSE_AHBIol0I
)
,
.CORETSE_AHBIiO1I
(
CORETSE_AHBo1i1I
)
,
.CORETSE_AHBliO1I
(
CORETSE_AHBiol1I
)
,
.CORETSE_AHBll0
(
CORETSE_AHBll0
)
,
.CORETSE_AHBoiO1I
(
CORETSE_AHBOOi1I
)
,
.CORETSE_AHBol0
(
CORETSE_AHBol0
)
,
.CORETSE_AHBil0
(
CORETSE_AHBil0
)
,
.CORETSE_AHBO00
(
CORETSE_AHBO00
)
,
.CORETSE_AHBI00
(
CORETSE_AHBI00
)
,
.CORETSE_AHBiiO1I
(
CORETSE_AHBIIi1I
)
,
.CORETSE_AHBIOI1I
(
CORETSE_AHBiio1I
)
,
.CORETSE_AHBoOI1I
(
CORETSE_AHBI1l1I
)
,
.CORETSE_AHBlOI1I
(
CORETSE_AHBiiI1I
)
,
.CORETSE_AHBOOI1I
(
CORETSE_AHBOli1I
)
)
;
endmodule
