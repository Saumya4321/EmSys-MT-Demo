// REVISION    : $Revision: 1.4 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
petbm
#
(
parameter
CORETSE_AHBlOI
=
1
'b
0
)
(
CORETSE_AHBi01
,
CORETSE_AHBO11
,
CORETSE_AHBI11
,
CORETSE_AHBl11
,
CORETSE_AHBl011
,
CORETSE_AHBl1O1
,
CORETSE_AHBo1O1
,
CORETSE_AHBi1O1
,
CORETSE_AHBOoO1
,
CORETSE_AHBIoO1
,
CORETSE_AHBloO1
,
CORETSE_AHBooO1
,
CORETSE_AHBooi0
,
CORETSE_AHBo01
,
CORETSE_AHBIo01
,
CORETSE_AHBlo01
,
CORETSE_AHBoo01
,
CORETSE_AHBiIO1
,
CORETSE_AHBOlO1
,
CORETSE_AHBio01
,
CORETSE_AHBIlO1
,
CORETSE_AHBOi01
,
CORETSE_AHBolO1
,
CORETSE_AHBIi01
,
CORETSE_AHBO0O1
,
CORETSE_AHBI0O1
,
CORETSE_AHBl0O1
,
CORETSE_AHBli01
,
CORETSE_AHBoi01
,
CORETSE_AHBo0O1
,
CORETSE_AHBii01
,
CORETSE_AHBi0O1
,
CORETSE_AHBO1O1
,
CORETSE_AHBOO11
,
CORETSE_AHBIO11
,
CORETSE_AHBoii0
,
CORETSE_AHBOOO1
,
CORETSE_AHBlO11
,
CORETSE_AHBoO11
,
CORETSE_AHBo011
)
;
input
CORETSE_AHBi01
;
input
CORETSE_AHBO11
;
input
CORETSE_AHBI11
;
input
CORETSE_AHBl11
;
input
CORETSE_AHBl011
;
input
CORETSE_AHBl1O1
;
input
CORETSE_AHBo1O1
;
input
CORETSE_AHBi1O1
;
input
[
15
:
0
]
CORETSE_AHBOoO1
;
input
[
15
:
0
]
CORETSE_AHBIoO1
;
input
CORETSE_AHBloO1
;
input
CORETSE_AHBooO1
;
input
[
4
:
0
]
CORETSE_AHBooi0
;
output
CORETSE_AHBo01
;
output
CORETSE_AHBIo01
;
output
CORETSE_AHBlo01
;
output
[
1
:
0
]
CORETSE_AHBoo01
;
output
CORETSE_AHBiIO1
;
output
CORETSE_AHBOlO1
;
output
CORETSE_AHBio01
;
output
[
15
:
0
]
CORETSE_AHBIlO1
;
output
CORETSE_AHBOi01
;
output
[
15
:
0
]
CORETSE_AHBolO1
;
output
CORETSE_AHBIi01
;
output
CORETSE_AHBO0O1
;
output
CORETSE_AHBI0O1
;
output
CORETSE_AHBl0O1
;
output
[
2
:
0
]
CORETSE_AHBli01
;
output
[
9
:
0
]
CORETSE_AHBoi01
;
output
CORETSE_AHBo0O1
;
output
CORETSE_AHBii01
;
output
CORETSE_AHBi0O1
;
output
CORETSE_AHBO1O1
;
output
CORETSE_AHBOO11
;
output
CORETSE_AHBIO11
;
output
CORETSE_AHBoii0
;
output
CORETSE_AHBOOO1
;
output
CORETSE_AHBlO11
;
output
CORETSE_AHBoO11
;
output
CORETSE_AHBo011
;
wire
CORETSE_AHBo01
;
reg
CORETSE_AHBIo01
;
reg
CORETSE_AHBlo01
;
reg
[
1
:
0
]
CORETSE_AHBoo01
;
reg
CORETSE_AHBiIO1
;
reg
CORETSE_AHBOlO1
;
reg
CORETSE_AHBio01
;
reg
[
15
:
0
]
CORETSE_AHBIlO1
;
reg
[
15
:
0
]
CORETSE_AHBolO1
;
wire
CORETSE_AHBOi01
;
wire
CORETSE_AHBIi01
;
reg
CORETSE_AHBO0O1
;
reg
CORETSE_AHBI0O1
;
reg
CORETSE_AHBl0O1
;
reg
[
2
:
0
]
CORETSE_AHBli01
;
reg
[
9
:
0
]
CORETSE_AHBoi01
;
reg
CORETSE_AHBo0O1
;
reg
CORETSE_AHBii01
;
reg
CORETSE_AHBi0O1
;
reg
CORETSE_AHBO1O1
;
reg
CORETSE_AHBOO11
;
reg
CORETSE_AHBIO11
;
reg
CORETSE_AHBoii0
;
reg
CORETSE_AHBOOO1
;
reg
CORETSE_AHBlO11
;
reg
CORETSE_AHBoO11
;
reg
CORETSE_AHBo011
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBilOII
;
wire
CORETSE_AHBO0OII
;
reg
CORETSE_AHBi1io
;
wire
[
5
:
0
]
CORETSE_AHBI0OII
;
reg
[
5
:
0
]
CORETSE_AHBl0OII
;
wire
CORETSE_AHBo0OII
;
reg
CORETSE_AHBi0OII
;
wire
CORETSE_AHBO1OII
;
reg
CORETSE_AHBI1OII
;
wire
CORETSE_AHBl1OII
;
wire
[
4
:
0
]
CORETSE_AHBo1OII
;
reg
[
4
:
0
]
CORETSE_AHBi1OII
;
wire
CORETSE_AHBOoOII
;
wire
[
4
:
0
]
CORETSE_AHBIoOII
;
reg
[
4
:
0
]
CORETSE_AHBloOII
;
wire
CORETSE_AHBooOII
;
reg
CORETSE_AHBioOII
;
wire
[
15
:
0
]
CORETSE_AHBOiOII
;
reg
[
15
:
0
]
CORETSE_AHBIiOII
;
reg
CORETSE_AHBliOII
,
CORETSE_AHBoiOII
,
CORETSE_AHBiiOII
;
reg
CORETSE_AHBOOIII
,
CORETSE_AHBIOIII
,
CORETSE_AHBlOIII
;
wire
[
15
:
0
]
CORETSE_AHBoOIII
,
CORETSE_AHBiOIII
;
reg
[
15
:
0
]
CORETSE_AHBOIIII
;
wire
CORETSE_AHBIIIII
,
CORETSE_AHBlIIII
,
CORETSE_AHBoIIII
,
CORETSE_AHBiIIII
,
CORETSE_AHBOlIII
;
wire
CORETSE_AHBIlIII
,
CORETSE_AHBllIII
,
CORETSE_AHBolIII
,
CORETSE_AHBilIII
,
CORETSE_AHBO0III
;
wire
CORETSE_AHBI0III
,
CORETSE_AHBl0III
,
CORETSE_AHBo0III
,
CORETSE_AHBi0III
,
CORETSE_AHBO1III
;
wire
CORETSE_AHBI1III
,
CORETSE_AHBl1III
,
CORETSE_AHBo1III
,
CORETSE_AHBi1III
,
CORETSE_AHBOoIII
;
wire
CORETSE_AHBIoIII
;
reg
CORETSE_AHBloIII
;
wire
CORETSE_AHBooIII
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBilOII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBilOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBO11
;
end
assign
CORETSE_AHBO0OII
=
~
CORETSE_AHBi1io
&
CORETSE_AHBI11
&
CORETSE_AHBO11
&
~
CORETSE_AHBilOII
|
CORETSE_AHBi1io
&
CORETSE_AHBI11
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBi1io
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBi1io
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0OII
;
end
assign
CORETSE_AHBI0OII
=
{
6
{
CORETSE_AHBi1io
&
CORETSE_AHBl0OII
<
6
'h
1e
}
}
&
CORETSE_AHBl0OII
+
6
'h
1
|
{
6
{
CORETSE_AHBioOII
&
CORETSE_AHBl0OII
<
6
'h
1e
}
}
&
CORETSE_AHBl0OII
+
6
'h
1
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBl0OII
[
5
:
0
]
<=
#
CORETSE_AHBIoII
6
'h
0
;
else
CORETSE_AHBl0OII
[
5
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0OII
[
5
:
0
]
;
end
assign
CORETSE_AHBo0OII
=
~
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
1
&
~
CORETSE_AHBO11
&
CORETSE_AHBilOII
|
CORETSE_AHBi0OII
&
CORETSE_AHBi1io
|
CORETSE_AHBi0OII
&
CORETSE_AHBioOII
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBi0OII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBi0OII
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0OII
;
end
assign
CORETSE_AHBO1OII
=
~
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1
&
CORETSE_AHBO11
&
~
CORETSE_AHBilOII
|
CORETSE_AHBI1OII
&
CORETSE_AHBI11
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBI1OII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBI1OII
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1OII
;
end
assign
CORETSE_AHBl1OII
=
(
CORETSE_AHBi0OII
|
CORETSE_AHBI1OII
)
&
CORETSE_AHBl0OII
[
5
:
0
]
>=
6
'h
2
&
CORETSE_AHBl0OII
[
5
:
0
]
<=
6
'h
6
;
assign
CORETSE_AHBo1OII
=
{
5
{
CORETSE_AHBl1OII
}
}
&
{
CORETSE_AHBi1OII
[
3
:
0
]
,
CORETSE_AHBO11
}
|
{
5
{
~
CORETSE_AHBl1OII
}
}
&
CORETSE_AHBi1OII
[
4
:
0
]
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBi1OII
[
4
:
0
]
<=
#
CORETSE_AHBIoII
5
'h
0
;
else
CORETSE_AHBi1OII
[
4
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1OII
[
4
:
0
]
;
end
assign
CORETSE_AHBOoOII
=
(
CORETSE_AHBi0OII
|
CORETSE_AHBI1OII
)
&
CORETSE_AHBl0OII
[
5
:
0
]
>=
6
'h
7
&
CORETSE_AHBl0OII
[
5
:
0
]
<=
6
'h
b
;
assign
CORETSE_AHBIoOII
=
{
5
{
CORETSE_AHBOoOII
}
}
&
{
CORETSE_AHBloOII
[
3
:
0
]
,
CORETSE_AHBO11
}
|
{
5
{
~
CORETSE_AHBOoOII
}
}
&
CORETSE_AHBloOII
[
4
:
0
]
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBloOII
[
4
:
0
]
<=
#
CORETSE_AHBIoII
5
'h
0
;
else
CORETSE_AHBloOII
[
4
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoOII
[
4
:
0
]
;
end
assign
CORETSE_AHBooOII
=
~
CORETSE_AHBioOII
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
c
&
~
CORETSE_AHBI11
|
CORETSE_AHBioOII
&
CORETSE_AHBl0OII
>
6
'h
c
&
CORETSE_AHBl0OII
<
6
'h
1e
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBioOII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBioOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBooOII
;
end
assign
CORETSE_AHBOiOII
=
{
16
{
CORETSE_AHBl0OII
>
6
'h
d
&
CORETSE_AHBI1OII
&
CORETSE_AHBI11
}
}
&
{
CORETSE_AHBIiOII
[
14
:
0
]
,
CORETSE_AHBO11
}
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBIiOII
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBIiOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiOII
;
end
assign
CORETSE_AHBoOIII
=
{
16
{
CORETSE_AHBI0III
}
}
&
{
CORETSE_AHBIo01
,
CORETSE_AHBlo01
,
CORETSE_AHBoo01
[
0
]
,
CORETSE_AHBiIO1
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBOlO1
,
CORETSE_AHBio01
,
1
'b
0
,
CORETSE_AHBoo01
[
1
]
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
,
1
'b
0
}
|
{
16
{
CORETSE_AHBl0III
}
}
&
{
4
'h
0
,
1
'h
0
,
1
'h
0
,
1
'h
0
,
1
'b
1
,
1
'h
0
,
1
'b
1
,
CORETSE_AHBl1O1
,
CORETSE_AHBo1O1
,
1
'b
1
,
CORETSE_AHBi1O1
,
1
'h
0
,
1
'b
1
}
|
{
16
{
CORETSE_AHBo0III
}
}
&
CORETSE_AHBIlO1
[
15
:
0
]
|
{
16
{
CORETSE_AHBi0III
}
}
&
CORETSE_AHBOoO1
[
15
:
0
]
|
{
16
{
CORETSE_AHBO1III
}
}
&
{
13
'h
0
,
1
'b
1
,
CORETSE_AHBloO1
,
1
'b
0
}
|
{
16
{
CORETSE_AHBI1III
}
}
&
CORETSE_AHBolO1
[
15
:
0
]
|
{
16
{
CORETSE_AHBl1III
}
}
&
CORETSE_AHBIoO1
[
15
:
0
]
|
{
16
{
CORETSE_AHBo1III
}
}
&
16
'h
a000
|
{
16
{
CORETSE_AHBi1III
}
}
&
{
CORETSE_AHBl0O1
,
CORETSE_AHBli01
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBoi01
}
|
{
16
{
CORETSE_AHBOoIII
}
}
&
{
CORETSE_AHBii01
,
CORETSE_AHBi0O1
,
CORETSE_AHBOO11
,
CORETSE_AHBIO11
,
CORETSE_AHBO1O1
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBo0O1
,
1
'b
0
,
CORETSE_AHBo011
,
CORETSE_AHBoO11
,
CORETSE_AHBlO11
,
1
'b
0
,
1
'b
0
,
CORETSE_AHBoii0
,
CORETSE_AHBOOO1
}
;
assign
CORETSE_AHBiOIII
=
{
16
{
CORETSE_AHBl0OII
==
6
'h
d
&
CORETSE_AHBioOII
}
}
&
{
CORETSE_AHBoOIII
[
15
:
0
]
}
|
{
16
{
CORETSE_AHBl0OII
>
6
'h
d
&
CORETSE_AHBioOII
}
}
&
{
CORETSE_AHBOIIII
[
14
:
0
]
,
1
'b
0
}
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBOIIII
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
CORETSE_AHBOIIII
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOIII
;
end
assign
CORETSE_AHBo01
=
(
(
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
)
&
CORETSE_AHBioOII
&
CORETSE_AHBl0OII
==
6
'h
d
)
&
CORETSE_AHBI11
|
(
(
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
)
&
CORETSE_AHBioOII
&
CORETSE_AHBl0OII
>
6
'h
d
)
&
CORETSE_AHBOIIII
[
15
]
|
~
(
(
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
)
&
CORETSE_AHBioOII
&
CORETSE_AHBl0OII
>=
6
'h
d
)
&
CORETSE_AHBl11
;
assign
CORETSE_AHBIIIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
00
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBI0III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
00
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBliOII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBliOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIIII
&
CORETSE_AHBIiOII
[
15
]
|
CORETSE_AHBliOII
&
~
CORETSE_AHBIo01
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
{
CORETSE_AHBlo01
,
CORETSE_AHBoo01
[
0
]
,
CORETSE_AHBiIO1
,
CORETSE_AHBio01
,
CORETSE_AHBoo01
[
1
]
}
<=
#
CORETSE_AHBIoII
5
'h
0
;
else
if
(
CORETSE_AHBIIIII
)
{
CORETSE_AHBlo01
,
CORETSE_AHBoo01
[
0
]
,
CORETSE_AHBiIO1
,
CORETSE_AHBio01
,
CORETSE_AHBoo01
[
1
]
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBIiOII
[
14
:
12
]
,
CORETSE_AHBIiOII
[
8
]
,
CORETSE_AHBIiOII
[
6
]
}
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBOOIII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOOIII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIIII
&
CORETSE_AHBIiOII
[
9
]
|
CORETSE_AHBOOIII
&
~
CORETSE_AHBOlO1
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBoiOII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBoiOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBliOII
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBiiOII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBiiOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBliOII
|
CORETSE_AHBoiOII
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBIo01
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBIo01
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiOII
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBIOIII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBIOIII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOIII
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBlOIII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBlOIII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOIII
|
CORETSE_AHBIOIII
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBOlO1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOlO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOIII
;
end
assign
CORETSE_AHBlIIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
01
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBl0III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
01
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBoIIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
04
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBo0III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
04
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBOi01
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
04
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBIlO1
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBoIIII
)
CORETSE_AHBIlO1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIiOII
;
end
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBI0O1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBIlIII
)
CORETSE_AHBI0O1
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBooO1
)
CORETSE_AHBI0O1
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
assign
CORETSE_AHBiIIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
05
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBi0III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
05
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBOlIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
06
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBO1III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
06
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBIoIII
=
CORETSE_AHBloO1
&
CORETSE_AHBO1III
|
CORETSE_AHBloIII
&
~
CORETSE_AHBO1III
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBloIII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBloIII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoIII
;
end
assign
CORETSE_AHBooIII
=
CORETSE_AHBloO1
&
CORETSE_AHBO1III
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBO0O1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO0O1
<=
#
CORETSE_AHBIoII
CORETSE_AHBooIII
;
end
assign
CORETSE_AHBIlIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
07
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBI1III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
07
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBIi01
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
07
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
CORETSE_AHBolO1
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBIlIII
)
CORETSE_AHBolO1
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIiOII
[
15
:
0
]
;
end
assign
CORETSE_AHBllIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
08
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBl1III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
08
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBolIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
0f
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBo1III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
0f
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
assign
CORETSE_AHBilIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
10
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBi1III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
10
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
{
CORETSE_AHBl0O1
,
CORETSE_AHBli01
,
CORETSE_AHBoi01
}
<=
#
CORETSE_AHBIoII
14
'h
0
;
else
if
(
CORETSE_AHBilIII
)
{
CORETSE_AHBl0O1
,
CORETSE_AHBli01
,
CORETSE_AHBoi01
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBIiOII
[
15
]
,
CORETSE_AHBIiOII
[
14
:
12
]
,
CORETSE_AHBIiOII
[
9
:
0
]
}
;
end
assign
CORETSE_AHBO0III
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
11
&
CORETSE_AHBI1OII
&
CORETSE_AHBl0OII
==
6
'h
1e
;
assign
CORETSE_AHBOoIII
=
CORETSE_AHBi1OII
[
4
:
0
]
==
CORETSE_AHBooi0
[
4
:
0
]
&
CORETSE_AHBloOII
[
4
:
0
]
==
5
'h
11
&
CORETSE_AHBi0OII
&
CORETSE_AHBl0OII
==
6
'h
d
;
always
@
(
posedge
CORETSE_AHBi01
or
posedge
CORETSE_AHBl011
)
begin
if
(
CORETSE_AHBl011
)
{
CORETSE_AHBii01
,
CORETSE_AHBi0O1
,
CORETSE_AHBOO11
,
CORETSE_AHBIO11
,
CORETSE_AHBO1O1
,
CORETSE_AHBo0O1
,
CORETSE_AHBo011
,
CORETSE_AHBoO11
,
CORETSE_AHBlO11
,
CORETSE_AHBoii0
,
CORETSE_AHBOOO1
}
<=
#
CORETSE_AHBIoII
11
'h
0
;
else
if
(
CORETSE_AHBO0III
)
{
CORETSE_AHBii01
,
CORETSE_AHBi0O1
,
CORETSE_AHBOO11
,
CORETSE_AHBIO11
,
CORETSE_AHBO1O1
,
CORETSE_AHBo0O1
,
CORETSE_AHBo011
,
CORETSE_AHBoO11
,
CORETSE_AHBlO11
,
CORETSE_AHBoii0
,
CORETSE_AHBOOO1
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBIiOII
[
15
:
12
]
,
CORETSE_AHBIiOII
[
11
]
,
CORETSE_AHBIiOII
[
8
]
,
CORETSE_AHBIiOII
[
6
:
4
]
,
CORETSE_AHBIiOII
[
1
:
0
]
}
;
end
endmodule
