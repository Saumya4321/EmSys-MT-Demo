// REVISION    : $Revision: 1.1 $
//         Mentor Graphics Corporation Proprietary and Confidential
//         Copyright Mentor Graphics Corporation and Licensors 2004
`timescale 1ps/1ps
module
arfque
(
CORETSE_AHBo0Ol
,
CORETSE_AHBi0Ol
,
CORETSE_AHBoio
,
CORETSE_AHBioo
,
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBO1Ol
,
CORETSE_AHBIlo
,
CORETSE_AHBI1Ol
,
CORETSE_AHBl1Ol
,
CORETSE_AHBo1Ol
,
CORETSE_AHBi1Ol
,
CORETSE_AHBOoOl
)
;
input
CORETSE_AHBo0Ol
;
input
CORETSE_AHBi0Ol
;
input
CORETSE_AHBoio
;
input
[
31
:
0
]
CORETSE_AHBioo
;
input
CORETSE_AHBOio
;
input
CORETSE_AHBIio
;
input
[
1
:
0
]
CORETSE_AHBlio
;
input
CORETSE_AHBO1Ol
;
output
CORETSE_AHBIlo
;
output
CORETSE_AHBI1Ol
;
output
[
31
:
0
]
CORETSE_AHBl1Ol
;
output
CORETSE_AHBo1Ol
;
output
CORETSE_AHBi1Ol
;
output
[
1
:
0
]
CORETSE_AHBOoOl
;
parameter
CORETSE_AHBIoII
=
1
;
reg
[
35
:
0
]
CORETSE_AHBIoOl
;
reg
[
35
:
0
]
CORETSE_AHBloOl
;
reg
[
1
:
0
]
CORETSE_AHBooOl
;
always
@
(
posedge
CORETSE_AHBo0Ol
or
negedge
CORETSE_AHBi0Ol
)
begin
if
(
~
CORETSE_AHBi0Ol
)
CORETSE_AHBIoOl
<=
#
CORETSE_AHBIoII
36
'h
0
;
else
if
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
)
CORETSE_AHBIoOl
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBioo
}
;
end
always
@
(
posedge
CORETSE_AHBo0Ol
or
negedge
CORETSE_AHBi0Ol
)
begin
if
(
~
CORETSE_AHBi0Ol
)
CORETSE_AHBooOl
[
0
]
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
)
&
~
(
CORETSE_AHBI1Ol
&
CORETSE_AHBO1Ol
)
&
CORETSE_AHBooOl
[
1
]
)
CORETSE_AHBooOl
[
0
]
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
~
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
)
&
(
CORETSE_AHBI1Ol
&
CORETSE_AHBO1Ol
)
)
CORETSE_AHBooOl
[
0
]
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBo0Ol
or
negedge
CORETSE_AHBi0Ol
)
begin
if
(
~
CORETSE_AHBi0Ol
)
CORETSE_AHBloOl
<=
#
CORETSE_AHBIoII
36
'h
0
;
else
if
(
(
CORETSE_AHBI1Ol
&
CORETSE_AHBO1Ol
)
&
CORETSE_AHBooOl
[
0
]
)
CORETSE_AHBloOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoOl
;
else
if
(
(
CORETSE_AHBI1Ol
&
CORETSE_AHBO1Ol
)
&
~
CORETSE_AHBooOl
[
0
]
)
CORETSE_AHBloOl
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBioo
}
;
else
if
(
~
CORETSE_AHBooOl
[
1
]
&
CORETSE_AHBooOl
[
0
]
)
CORETSE_AHBloOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoOl
;
else
if
(
~
CORETSE_AHBooOl
[
1
]
&
~
CORETSE_AHBooOl
[
0
]
)
CORETSE_AHBloOl
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBioo
}
;
end
always
@
(
posedge
CORETSE_AHBo0Ol
or
negedge
CORETSE_AHBi0Ol
)
begin
if
(
~
CORETSE_AHBi0Ol
)
CORETSE_AHBooOl
[
1
]
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBooOl
[
0
]
|
(
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
)
&
~
(
CORETSE_AHBI1Ol
&
CORETSE_AHBO1Ol
)
)
)
CORETSE_AHBooOl
[
1
]
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
(
~
(
CORETSE_AHBoio
&
CORETSE_AHBIlo
)
&
(
CORETSE_AHBI1Ol
&
CORETSE_AHBO1Ol
)
)
)
CORETSE_AHBooOl
[
1
]
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
assign
{
CORETSE_AHBo1Ol
,
CORETSE_AHBi1Ol
,
CORETSE_AHBOoOl
,
CORETSE_AHBl1Ol
}
=
CORETSE_AHBloOl
;
assign
CORETSE_AHBI1Ol
=
CORETSE_AHBooOl
[
1
]
;
assign
CORETSE_AHBIlo
=
~
CORETSE_AHBooOl
[
0
]
;
endmodule
