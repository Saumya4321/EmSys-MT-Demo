// REVISION    : $Revision: 1.1 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_cnvrxo
(
CORETSE_AHBOI10
,
CORETSE_AHBii0
,
CORETSE_AHBo11
,
CORETSE_AHBOo10
,
CORETSE_AHBIo10
,
CORETSE_AHBlo10
,
CORETSE_AHBoo10
,
CORETSE_AHBio10
,
CORETSE_AHBlI
,
CORETSE_AHBiI
,
CORETSE_AHBIl
,
CORETSE_AHBi110
)
;
input
CORETSE_AHBOI10
;
input
CORETSE_AHBii0
;
input
[
1
:
0
]
CORETSE_AHBo11
;
input
[
7
:
0
]
CORETSE_AHBOo10
;
input
CORETSE_AHBIo10
;
input
CORETSE_AHBlo10
;
input
CORETSE_AHBoo10
;
input
[
3
:
0
]
CORETSE_AHBio10
;
output
[
7
:
0
]
CORETSE_AHBlI
;
output
CORETSE_AHBiI
;
output
CORETSE_AHBIl
;
output
[
3
:
0
]
CORETSE_AHBi110
;
`define CORETSE_AHBIoII  \
# \
1
reg
[
7
:
0
]
CORETSE_AHBlI
;
reg
CORETSE_AHBiI
;
reg
CORETSE_AHBIl
;
reg
[
3
:
0
]
CORETSE_AHBi110
;
reg
CORETSE_AHBo1o0
;
reg
[
2
:
0
]
CORETSE_AHBI1o0
;
wire
CORETSE_AHBi1o0
;
wire
[
7
:
0
]
CORETSE_AHBOoo0
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBOI10
)
begin
if
(
CORETSE_AHBOI10
)
CORETSE_AHBI1o0
<=
`CORETSE_AHBIoII
3
'h
0
;
else
CORETSE_AHBI1o0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBI1o0
[
1
:
0
]
,
CORETSE_AHBoo10
}
;
end
assign
CORETSE_AHBi1o0
=
CORETSE_AHBI1o0
[
1
]
&
~
CORETSE_AHBI1o0
[
2
]
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBOI10
)
begin
if
(
CORETSE_AHBOI10
)
CORETSE_AHBo1o0
<=
`CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1o0
&
~
CORETSE_AHBIo10
)
CORETSE_AHBo1o0
<=
`CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBo1o0
<=
`CORETSE_AHBIoII
~
CORETSE_AHBo1o0
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBOI10
)
begin
if
(
CORETSE_AHBOI10
)
CORETSE_AHBi110
<=
`CORETSE_AHBIoII
4
'h
4
;
else
if
(
(
CORETSE_AHBo11
==
2
'b
10
)
&
CORETSE_AHBi1o0
&
~
CORETSE_AHBIo10
)
CORETSE_AHBi110
<=
`CORETSE_AHBIoII
{
CORETSE_AHBio10
[
2
:
0
]
,
1
'b
0
}
;
else
if
(
(
CORETSE_AHBo11
!=
2
'b
10
)
&
CORETSE_AHBi1o0
&
~
CORETSE_AHBIo10
)
CORETSE_AHBi110
<=
`CORETSE_AHBIoII
CORETSE_AHBio10
;
else
if
(
(
~
CORETSE_AHBo1o0
)
|
(
CORETSE_AHBo11
==
2
'b
10
)
)
CORETSE_AHBi110
<=
`CORETSE_AHBIoII
CORETSE_AHBi110
+
4
'h
1
;
end
assign
CORETSE_AHBOoo0
=
{
8
{
(
CORETSE_AHBo11
==
2
'h
2
)
}
}
&
CORETSE_AHBOo10
|
{
8
{
(
CORETSE_AHBo11
!=
2
'h
2
)
&
CORETSE_AHBo1o0
}
}
&
{
4
'h
0
,
CORETSE_AHBOo10
[
3
:
0
]
}
|
{
8
{
(
CORETSE_AHBo11
!=
2
'h
2
)
&
~
CORETSE_AHBo1o0
}
}
&
{
4
'h
0
,
CORETSE_AHBOo10
[
7
:
4
]
}
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBOI10
)
begin
if
(
CORETSE_AHBOI10
)
CORETSE_AHBlI
<=
`CORETSE_AHBIoII
8
'h
0
;
else
CORETSE_AHBlI
<=
`CORETSE_AHBIoII
CORETSE_AHBOoo0
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBOI10
)
begin
if
(
CORETSE_AHBOI10
)
CORETSE_AHBiI
<=
`CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiI
<=
`CORETSE_AHBIoII
CORETSE_AHBIo10
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBOI10
)
begin
if
(
CORETSE_AHBOI10
)
CORETSE_AHBIl
<=
`CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIl
<=
`CORETSE_AHBIoII
CORETSE_AHBlo10
;
end
endmodule
