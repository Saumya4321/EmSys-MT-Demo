// REVISION    : $Revision: 1.1 $
//              Mentor Proprietary and Confidential
//              Copyright (c) 2000, Mentor Intellectual Property Development
`timescale 1ns/1ns
module
pemstat_store
(
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
,
CORETSE_AHBiOIi
,
CORETSE_AHBOIIi
,
CORETSE_AHBIIIi
,
CORETSE_AHBlIIi
,
CORETSE_AHBoIIi
,
CORETSE_AHBiIIi
,
CORETSE_AHBl1li
,
CORETSE_AHBOlIi
,
CORETSE_AHBIlIi
,
CORETSE_AHBllIi
,
CORETSE_AHBolIi
,
CORETSE_AHBilIi
,
CORETSE_AHBO0Ii
,
CORETSE_AHBI0Ii
,
CORETSE_AHBl0Ii
,
CORETSE_AHBo0Ii
,
CORETSE_AHBi0Ii
,
CORETSE_AHBO1Ii
,
CORETSE_AHBI1Ii
,
CORETSE_AHBl1Ii
,
CORETSE_AHBo1Ii
,
CORETSE_AHBi1Ii
,
CORETSE_AHBOoIi
,
CORETSE_AHBIoIi
,
CORETSE_AHBloIi
,
CORETSE_AHBooIi
,
CORETSE_AHBioIi
,
CORETSE_AHBOiIi
,
CORETSE_AHBIiIi
,
CORETSE_AHBliIi
,
CORETSE_AHBoiIi
,
CORETSE_AHBiiIi
,
CORETSE_AHBOOli
,
CORETSE_AHBIOli
,
CORETSE_AHBlOli
,
CORETSE_AHBoOli
,
CORETSE_AHBiOli
,
CORETSE_AHBOIli
,
CORETSE_AHBIIli
,
CORETSE_AHBlIli
,
CORETSE_AHBoIli
,
CORETSE_AHBiIli
,
CORETSE_AHBOlli
,
CORETSE_AHBIlli
,
CORETSE_AHBllli
,
CORETSE_AHBolli
,
CORETSE_AHBilli
,
CORETSE_AHBO0li
,
CORETSE_AHBI0li
,
CORETSE_AHBl0li
,
CORETSE_AHBo0li
,
CORETSE_AHBi0li
)
;
input
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
;
input
[
15
:
0
]
CORETSE_AHBiOIi
;
input
[
3
:
0
]
CORETSE_AHBOIIi
;
input
[
43
:
0
]
CORETSE_AHBIIIi
;
input
[
43
:
0
]
CORETSE_AHBlIIi
;
input
[
43
:
0
]
CORETSE_AHBoIIi
;
input
[
43
:
0
]
CORETSE_AHBiIIi
;
input
[
31
:
0
]
CORETSE_AHBl1li
;
output
[
43
:
0
]
CORETSE_AHBOlIi
;
output
[
30
:
0
]
CORETSE_AHBIlIi
,
CORETSE_AHBllIi
,
CORETSE_AHBolIi
,
CORETSE_AHBilIi
,
CORETSE_AHBO0Ii
,
CORETSE_AHBI0Ii
,
CORETSE_AHBl0Ii
,
CORETSE_AHBo0Ii
;
output
[
30
:
0
]
CORETSE_AHBi0Ii
,
CORETSE_AHBO1Ii
,
CORETSE_AHBI1Ii
,
CORETSE_AHBl1Ii
,
CORETSE_AHBo1Ii
,
CORETSE_AHBi1Ii
,
CORETSE_AHBOoIi
,
CORETSE_AHBIoIi
;
output
[
30
:
0
]
CORETSE_AHBloIi
,
CORETSE_AHBooIi
,
CORETSE_AHBioIi
,
CORETSE_AHBOiIi
,
CORETSE_AHBIiIi
,
CORETSE_AHBliIi
,
CORETSE_AHBoiIi
,
CORETSE_AHBiiIi
;
output
[
30
:
0
]
CORETSE_AHBOOli
,
CORETSE_AHBIOli
,
CORETSE_AHBlOli
,
CORETSE_AHBoOli
,
CORETSE_AHBiOli
,
CORETSE_AHBOIli
,
CORETSE_AHBIIli
,
CORETSE_AHBlIli
;
output
[
30
:
0
]
CORETSE_AHBoIli
,
CORETSE_AHBiIli
,
CORETSE_AHBOlli
,
CORETSE_AHBIlli
,
CORETSE_AHBllli
,
CORETSE_AHBolli
,
CORETSE_AHBilli
,
CORETSE_AHBO0li
;
output
[
30
:
0
]
CORETSE_AHBI0li
,
CORETSE_AHBl0li
,
CORETSE_AHBo0li
,
CORETSE_AHBi0li
;
pemstat_linc
CORETSE_AHBOi0i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
00
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
00
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
00
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
00
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBIlIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
00
]
)
)
;
pemstat_linc
CORETSE_AHBIi0i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
01
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
01
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
01
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
01
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBllIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
01
]
)
)
;
pemstat_linc
CORETSE_AHBli0i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
02
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
02
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
02
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
02
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBolIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
02
]
)
)
;
pemstat_linc
CORETSE_AHBoi0i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
03
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
03
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
03
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
03
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBilIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
03
]
)
)
;
pemstat_linc
CORETSE_AHBii0i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
04
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
04
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
04
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
04
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBO0Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
04
]
)
)
;
pemstat_linc
CORETSE_AHBOO1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
05
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
05
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
05
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
05
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBI0Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
05
]
)
)
;
pemstat_linc
CORETSE_AHBIO1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
06
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
06
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
06
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
06
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBl0Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
06
]
)
)
;
pemstat_ladd
CORETSE_AHBlO1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBi10i
(
CORETSE_AHBIIIi
[
07
]
)
,
.CORETSE_AHBOo0i
(
CORETSE_AHBiOIi
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
07
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
07
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
07
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBo0Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
07
]
)
)
;
pemstat_linc
CORETSE_AHBoO1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
08
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
08
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
08
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
08
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBi0Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
08
]
)
)
;
pemstat_sinc
CORETSE_AHBiO1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
09
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
09
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
09
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
09
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBO1Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
09
]
)
)
;
pemstat_linc
CORETSE_AHBOI1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
10
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
10
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
10
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
10
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBI1Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
10
]
)
)
;
pemstat_linc
CORETSE_AHBII1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
11
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
11
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
11
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
11
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBl1Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
11
]
)
)
;
pemstat_sinc
CORETSE_AHBlI1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
12
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
12
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
12
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
12
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBo1Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
12
]
)
)
;
pemstat_sinc
CORETSE_AHBoI1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
13
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
13
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
13
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
13
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBi1Ii
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
13
]
)
)
;
pemstat_sinc
CORETSE_AHBiI1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
14
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
14
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
14
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
14
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBOoIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
14
]
)
)
;
pemstat_sinc
CORETSE_AHBOl1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
15
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
15
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
15
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
15
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBIoIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
15
]
)
)
;
pemstat_sinc
CORETSE_AHBIl1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
16
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
16
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
16
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
16
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBloIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
16
]
)
)
;
pemstat_sinc
CORETSE_AHBll1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
17
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
17
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
17
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
17
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBooIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
17
]
)
)
;
pemstat_sinc
CORETSE_AHBol1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
18
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
18
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
18
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
18
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBioIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
18
]
)
)
;
pemstat_sinc
CORETSE_AHBil1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
19
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
19
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
19
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
19
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBOiIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
19
]
)
)
;
pemstat_sinc
CORETSE_AHBO01i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
20
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
20
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
20
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
20
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBIiIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
20
]
)
)
;
pemstat_sinc
CORETSE_AHBI01i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
21
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
21
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
21
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
21
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBliIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
21
]
)
)
;
pemstat_sinc
CORETSE_AHBl01i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
22
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
22
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
22
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
22
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBoiIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
22
]
)
)
;
pemstat_sinc
CORETSE_AHBo01i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
23
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
23
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
23
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
23
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBiiIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
23
]
)
)
;
pemstat_ladd
CORETSE_AHBi01i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBi10i
(
CORETSE_AHBIIIi
[
24
]
)
,
.CORETSE_AHBOo0i
(
CORETSE_AHBiOIi
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
24
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
24
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
24
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBOOli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
24
]
)
)
;
pemstat_linc
CORETSE_AHBO11i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
25
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
25
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
25
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
25
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBIOli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
25
]
)
)
;
pemstat_linc
CORETSE_AHBI11i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
26
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
26
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
26
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
26
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBlOli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
26
]
)
)
;
pemstat_linc
CORETSE_AHBl11i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
27
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
27
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
27
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
27
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBoOli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
27
]
)
)
;
pemstat_sinc
CORETSE_AHBo11i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
28
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
28
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
28
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
28
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBiOli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
28
]
)
)
;
pemstat_sinchd
CORETSE_AHBi11i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
29
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
29
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
29
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
29
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBOIli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
29
]
)
)
;
pemstat_sinchd
CORETSE_AHBOo1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
30
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
30
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
30
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
30
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBIIli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
30
]
)
)
;
pemstat_sinchd
CORETSE_AHBIo1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
31
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
31
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
31
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
31
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBlIli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
31
]
)
)
;
pemstat_sinchd
CORETSE_AHBlo1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
32
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
32
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
32
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
32
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBoIli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
32
]
)
)
;
pemstat_sinchd
CORETSE_AHBoo1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
33
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
33
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
33
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
33
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBiIli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
33
]
)
)
;
pemstat_sinchd
CORETSE_AHBio1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
34
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
34
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
34
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
34
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBOlli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
34
]
)
)
;
pemstat_sadd
CORETSE_AHBOi1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBi10i
(
CORETSE_AHBIIIi
[
35
]
)
,
.CORETSE_AHBOo0i
(
CORETSE_AHBOIIi
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
35
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
35
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
35
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBIlli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
35
]
)
)
;
pemstat_sinc
CORETSE_AHBIi1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
36
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
36
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
36
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
36
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBllli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
36
]
)
)
;
pemstat_sinc
CORETSE_AHBli1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
37
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
37
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
37
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
37
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBolli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
37
]
)
)
;
pemstat_sincnf
CORETSE_AHBoi1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
38
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
38
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
38
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
38
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBilli
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
38
]
)
)
;
pemstat_sincnf
CORETSE_AHBii1i
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
39
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
39
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
39
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
39
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBO0li
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
39
]
)
)
;
pemstat_sincnf
CORETSE_AHBOOoi
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
40
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
40
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
40
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
40
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBI0li
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
40
]
)
)
;
pemstat_sincnf
CORETSE_AHBIOoi
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
41
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
41
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
41
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
41
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBl0li
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
41
]
)
)
;
pemstat_sincnf
CORETSE_AHBlOoi
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
42
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
42
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
42
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
42
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBo0li
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
42
]
)
)
;
pemstat_sincnf
CORETSE_AHBoOoi
(
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBio0i
(
CORETSE_AHBIIIi
[
43
]
)
,
.CORETSE_AHBoIIi
(
CORETSE_AHBoIIi
[
43
]
)
,
.CORETSE_AHBl1li
(
CORETSE_AHBl1li
[
30
:
0
]
)
,
.CORETSE_AHBiIIi
(
CORETSE_AHBiIIi
[
43
]
)
,
.CORETSE_AHBlIIi
(
CORETSE_AHBlIIi
[
43
]
)
,
.CORETSE_AHBIo0i
(
CORETSE_AHBi0li
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBOlIi
[
43
]
)
)
;
endmodule
