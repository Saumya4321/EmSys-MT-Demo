//                        Proprietary and Confidential 
// REVISION    : $Revision: $ 
`include "include.v"
module
ptp_hstinf
#
(
parameter
CORETSE_AHBlII
=
2
,
parameter
CORETSE_AHBIII
=
1
,
parameter
CORETSE_AHBiII
=
2
,
parameter
CORETSE_AHBoII
=
1
,
parameter
CORETSE_AHBOlI
=
18
,
parameter
CORETSE_AHBIlI
=
18
,
parameter
CORETSE_AHBllI
=
5
,
parameter
CORETSE_AHBolI
=
5
)
(
input
CORETSE_AHBiil0,
input
CORETSE_AHBi10lI,
input
CORETSE_AHBOl0,
input
CORETSE_AHBOo0lI,
input
CORETSE_AHBIo0lI,
input
CORETSE_AHBlo0lI,
input
CORETSE_AHBoo0lI,
input
[
4
:
0
]
CORETSE_AHBoO00,
input
[
31
:
0
]
CORETSE_AHBio0lI,
input
[
79
:
0
]
CORETSE_AHBOi0lI,
input
CORETSE_AHBIi0lI,
input
CORETSE_AHBli0lI,
input
CORETSE_AHBoi0lI,
input
CORETSE_AHBii0lI,
input
CORETSE_AHBOO1lI,
input
[
3
:
0
]
CORETSE_AHBIO1lI,
input
[
15
:
0
]
CORETSE_AHBlO1lI,
input
[
79
:
0
]
CORETSE_AHBoO1lI,
input
[
79
:
0
]
CORETSE_AHBioo1,
input
[
3
:
0
]
CORETSE_AHBiO1lI,
input
[
15
:
0
]
CORETSE_AHBOI1lI,
input
[
79
:
0
]
CORETSE_AHBII1lI,
input
[
79
:
0
]
CORETSE_AHBlI1lI,
input
CORETSE_AHBlI0,
input
CORETSE_AHBoI0,
input
CORETSE_AHBiI0,
output
[
31
:
0
]
CORETSE_AHBoI1lI,
output
CORETSE_AHBiI1lI,
output
CORETSE_AHBOl1lI,
output
CORETSE_AHBIl1lI,
output
[
79
:
0
]
CORETSE_AHBll1lI,
output
[
79
:
0
]
CORETSE_AHBol1lI,
output
[
79
:
0
]
CORETSE_AHBil1lI,
output
[
7
:
0
]
CORETSE_AHBO01lI,
output
[
7
:
0
]
CORETSE_AHBI01lI,
output
CORETSE_AHBl01lI,
output
CORETSE_AHBo01lI,
output
CORETSE_AHBi01lI,
output
CORETSE_AHBO11lI,
output
CORETSE_AHBI11lI,
output
CORETSE_AHBl11lI,
output
CORETSE_AHBo11lI,
output
CORETSE_AHBi11lI,
output
[
`CORETSE_AHBIoI0
:
0
]
CORETSE_AHBOo1lI,
output
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
CORETSE_AHBIo1lI,
output
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
CORETSE_AHBlo1lI,
output
CORETSE_AHBoo1lI,
output
CORETSE_AHBio1lI,
output
CORETSE_AHBOi1lI,
output
CORETSE_AHBIi1lI,
output
CORETSE_AHBli1lI,
output
CORETSE_AHBoi1lI,
output
CORETSE_AHBii1lI
)
;
localparam
[
CORETSE_AHBllI
-
1
:
0
]
CORETSE_AHBOOolI
=
CORETSE_AHBOlI
;
localparam
[
CORETSE_AHBolI
-
1
:
0
]
CORETSE_AHBIOolI
=
CORETSE_AHBIlI
;
localparam
[
CORETSE_AHBllI
-
1
:
0
]
CORETSE_AHBlOolI
=
(
(
(
2
**
CORETSE_AHBllI
)
%
6
)
==
0
)
?
(
2
**
CORETSE_AHBllI
-
1
)
:
(
(
2
**
CORETSE_AHBllI
-
1
)
-
(
(
2
**
CORETSE_AHBllI
)
%
6
)
)
;
localparam
[
CORETSE_AHBolI
-
1
:
0
]
CORETSE_AHBoOolI
=
(
(
(
2
**
CORETSE_AHBolI
)
%
6
)
==
0
)
?
(
2
**
CORETSE_AHBolI
-
1
)
:
(
(
2
**
CORETSE_AHBolI
-
1
)
-
(
(
2
**
CORETSE_AHBolI
)
%
6
)
)
;
reg
[
31
:
0
]
CORETSE_AHBiOolI
;
wire
[
31
:
0
]
CORETSE_AHBOIolI
;
reg
[
31
:
0
]
CORETSE_AHBIIolI
;
wire
[
31
:
0
]
CORETSE_AHBlIolI
;
reg
[
15
:
0
]
CORETSE_AHBoIolI
;
wire
[
15
:
0
]
CORETSE_AHBiIolI
;
reg
[
31
:
0
]
CORETSE_AHBOlolI
;
wire
[
31
:
0
]
CORETSE_AHBIlolI
;
reg
[
31
:
0
]
CORETSE_AHBllolI
;
wire
[
31
:
0
]
CORETSE_AHBololI
;
reg
[
15
:
0
]
CORETSE_AHBilolI
;
wire
[
15
:
0
]
CORETSE_AHBO0olI
;
reg
[
31
:
0
]
CORETSE_AHBI0olI
;
wire
[
31
:
0
]
CORETSE_AHBl0olI
;
reg
[
31
:
0
]
CORETSE_AHBo0olI
;
wire
[
31
:
0
]
CORETSE_AHBi0olI
;
reg
[
15
:
0
]
CORETSE_AHBO1olI
;
wire
[
15
:
0
]
CORETSE_AHBI1olI
;
reg
[
31
:
0
]
CORETSE_AHBl1olI
;
wire
[
31
:
0
]
CORETSE_AHBo1olI
;
reg
[
31
:
0
]
CORETSE_AHBi1olI
;
wire
[
31
:
0
]
CORETSE_AHBOoolI
;
reg
[
15
:
0
]
CORETSE_AHBIoolI
;
wire
[
15
:
0
]
CORETSE_AHBloolI
;
reg
[
31
:
0
]
CORETSE_AHBooolI
;
wire
[
31
:
0
]
CORETSE_AHBioolI
;
reg
[
31
:
0
]
CORETSE_AHBOiolI
;
wire
[
31
:
0
]
CORETSE_AHBIiolI
;
reg
[
15
:
0
]
CORETSE_AHBliolI
;
wire
[
15
:
0
]
CORETSE_AHBoiolI
;
reg
[
7
:
0
]
CORETSE_AHBiiolI
;
wire
[
7
:
0
]
CORETSE_AHBOOilI
;
reg
[
7
:
0
]
CORETSE_AHBIOilI
;
wire
[
7
:
0
]
CORETSE_AHBlOilI
;
reg
CORETSE_AHBoOilI
;
wire
CORETSE_AHBiOilI
;
reg
[
`CORETSE_AHBO1I0
:
0
]
CORETSE_AHBOIilI
;
wire
[
`CORETSE_AHBO1I0
:
0
]
CORETSE_AHBIIilI
;
reg
[
9
:
0
]
CORETSE_AHBlIilI
;
wire
[
9
:
0
]
CORETSE_AHBoIilI
;
reg
[
10
:
0
]
CORETSE_AHBiIilI
;
wire
[
10
:
0
]
CORETSE_AHBOlilI
;
reg
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
CORETSE_AHBIlilI
;
wire
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
CORETSE_AHBllilI
;
reg
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
CORETSE_AHBolilI
;
wire
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
CORETSE_AHBililI
;
wire
CORETSE_AHBO0ilI
;
wire
CORETSE_AHBI0ilI
;
wire
CORETSE_AHBl0ilI
;
wire
CORETSE_AHBo0ilI
;
wire
CORETSE_AHBi0ilI
;
wire
CORETSE_AHBO1ilI
;
wire
CORETSE_AHBI1ilI
;
wire
CORETSE_AHBl1ilI
;
wire
CORETSE_AHBo1ilI
;
wire
CORETSE_AHBi1ilI
;
reg
CORETSE_AHBOoilI
;
wire
CORETSE_AHBIoilI
;
reg
CORETSE_AHBloilI
;
wire
CORETSE_AHBooilI
;
reg
CORETSE_AHBioilI
;
wire
CORETSE_AHBOiilI
;
reg
CORETSE_AHBIiilI
;
wire
CORETSE_AHBliilI
;
reg
CORETSE_AHBoiilI
;
wire
CORETSE_AHBiiilI
;
reg
CORETSE_AHBOOO0I
;
wire
CORETSE_AHBIOO0I
;
reg
CORETSE_AHBlOO0I
;
wire
CORETSE_AHBoOO0I
;
reg
[
5
:
0
]
CORETSE_AHBiOO0I
;
wire
[
5
:
0
]
CORETSE_AHBOIO0I
;
reg
CORETSE_AHBIIO0I
;
wire
CORETSE_AHBlIO0I
;
reg
CORETSE_AHBoIO0I
;
wire
CORETSE_AHBiIO0I
;
reg
CORETSE_AHBOlO0I
;
wire
CORETSE_AHBIlO0I
;
reg
CORETSE_AHBllO0I
;
wire
CORETSE_AHBolO0I
;
reg
CORETSE_AHBilO0I
;
wire
CORETSE_AHBO0O0I
;
reg
CORETSE_AHBI0O0I
;
wire
CORETSE_AHBl0O0I
;
reg
CORETSE_AHBo0O0I
;
wire
CORETSE_AHBi0O0I
;
reg
[
5
:
0
]
CORETSE_AHBO1O0I
;
wire
[
5
:
0
]
CORETSE_AHBI1O0I
;
wire
[
31
:
0
]
CORETSE_AHBl1O0I
;
wire
[
31
:
0
]
CORETSE_AHBo1O0I
;
wire
[
31
:
0
]
CORETSE_AHBi1O0I
;
wire
[
31
:
0
]
CORETSE_AHBOoO0I
;
wire
CORETSE_AHBIoO0I
;
wire
CORETSE_AHBloO0I
;
wire
CORETSE_AHBooO0I
;
wire
CORETSE_AHBioO0I
;
wire
CORETSE_AHBOiO0I
;
wire
CORETSE_AHBIiO0I
;
wire
CORETSE_AHBliO0I
;
wire
CORETSE_AHBoiO0I
;
reg
CORETSE_AHBiiO0I
;
reg
CORETSE_AHBOOI0I
;
reg
CORETSE_AHBIOI0I
;
reg
CORETSE_AHBlOI0I
;
reg
CORETSE_AHBoOI0I
;
reg
CORETSE_AHBiOI0I
;
wire
CORETSE_AHBOII0I
;
wire
CORETSE_AHBIII0I
;
reg
CORETSE_AHBlII0I
;
wire
CORETSE_AHBoII0I
;
wire
[
31
:
0
]
CORETSE_AHBiII0I
;
wire
CORETSE_AHBOlI0I
;
wire
CORETSE_AHBIlI0I
;
wire
CORETSE_AHBllI0I
;
wire
CORETSE_AHBolI0I
;
reg
CORETSE_AHBilI0I
;
reg
CORETSE_AHBO0I0I
;
reg
CORETSE_AHBI0I0I
;
wire
CORETSE_AHBl0I0I
;
reg
[
15
:
0
]
CORETSE_AHBo0I0I
;
wire
[
15
:
0
]
CORETSE_AHBi0I0I
;
reg
[
3
:
0
]
CORETSE_AHBO1I0I
;
wire
[
3
:
0
]
CORETSE_AHBI1I0I
;
reg
[
79
:
0
]
CORETSE_AHBl1I0I
;
wire
[
79
:
0
]
CORETSE_AHBo1I0I
;
reg
[
79
:
0
]
CORETSE_AHBi1I0I
;
wire
[
79
:
0
]
CORETSE_AHBOoI0I
;
reg
CORETSE_AHBIoI0I
;
reg
CORETSE_AHBloI0I
;
reg
CORETSE_AHBooI0I
;
reg
[
15
:
0
]
CORETSE_AHBioI0I
;
wire
[
15
:
0
]
CORETSE_AHBOiI0I
;
reg
[
3
:
0
]
CORETSE_AHBIiI0I
;
wire
[
3
:
0
]
CORETSE_AHBliI0I
;
reg
[
79
:
0
]
CORETSE_AHBoiI0I
;
wire
[
79
:
0
]
CORETSE_AHBiiI0I
;
reg
[
79
:
0
]
CORETSE_AHBOOl0I
;
wire
[
79
:
0
]
CORETSE_AHBIOl0I
;
wire
CORETSE_AHBlOl0I
;
wire
CORETSE_AHBoOl0I
;
wire
CORETSE_AHBiOl0I
;
wire
CORETSE_AHBOIl0I
;
wire
CORETSE_AHBIIl0I
;
reg
CORETSE_AHBlIl0I
;
reg
CORETSE_AHBoIl0I
;
reg
CORETSE_AHBiIl0I
;
reg
CORETSE_AHBOll0I
;
reg
CORETSE_AHBIll0I
;
wire
CORETSE_AHBlll0I
;
wire
CORETSE_AHBoll0I
,
CORETSE_AHBill0I
;
wire
CORETSE_AHBO0l0I
,
CORETSE_AHBI0l0I
;
wire
CORETSE_AHBl0l0I
,
CORETSE_AHBo0l0I
;
wire
CORETSE_AHBi0l0I
;
wire
CORETSE_AHBO1l0I
;
wire
CORETSE_AHBI1l0I
;
wire
CORETSE_AHBl1l0I
;
wire
CORETSE_AHBo1l0I
;
wire
CORETSE_AHBi1l0I
;
wire
CORETSE_AHBOol0I
;
reg
[
`CORETSE_AHBIoI0
:
0
]
CORETSE_AHBIol0I
;
wire
[
`CORETSE_AHBIoI0
:
0
]
CORETSE_AHBlol0I
;
reg
[
31
:
0
]
CORETSE_AHBool0I
;
wire
[
31
:
0
]
CORETSE_AHBiol0I
;
reg
[
31
:
0
]
CORETSE_AHBOil0I
;
wire
[
31
:
0
]
CORETSE_AHBIil0I
;
reg
[
31
:
0
]
CORETSE_AHBlil0I
;
wire
[
31
:
0
]
CORETSE_AHBoil0I
;
reg
[
31
:
0
]
CORETSE_AHBiil0I
;
wire
[
31
:
0
]
CORETSE_AHBOO00I
;
reg
[
31
:
0
]
CORETSE_AHBIO00I
;
wire
[
31
:
0
]
CORETSE_AHBlO00I
;
reg
[
31
:
0
]
CORETSE_AHBoO00I
;
wire
[
31
:
0
]
CORETSE_AHBiO00I
;
wire
CORETSE_AHBOI00I
;
wire
CORETSE_AHBII00I
;
wire
CORETSE_AHBlI00I
;
reg
CORETSE_AHBoI00I
;
reg
CORETSE_AHBiI00I
;
reg
CORETSE_AHBOl00I
;
reg
CORETSE_AHBIl00I
;
reg
CORETSE_AHBll00I
;
reg
CORETSE_AHBol00I
;
reg
CORETSE_AHBil00I
;
reg
CORETSE_AHBO000I
;
reg
CORETSE_AHBI000I
;
wire
CORETSE_AHBl000I
;
reg
CORETSE_AHBo000I
;
wire
CORETSE_AHBi000I
;
reg
CORETSE_AHBO100I
;
wire
CORETSE_AHBI100I
;
reg
CORETSE_AHBl100I
;
reg
CORETSE_AHBo100I
;
reg
CORETSE_AHBi100I
;
reg
CORETSE_AHBOo00I
;
reg
CORETSE_AHBIo00I
;
reg
CORETSE_AHBlo00I
;
reg
CORETSE_AHBoo00I
;
reg
CORETSE_AHBio00I
;
reg
CORETSE_AHBOi00I
;
reg
CORETSE_AHBIi00I
;
reg
CORETSE_AHBli00I
;
reg
CORETSE_AHBoi00I
;
reg
CORETSE_AHBii00I
;
reg
CORETSE_AHBOO10I
;
reg
CORETSE_AHBIO10I
;
reg
CORETSE_AHBlO10I
;
wire
CORETSE_AHBoO10I
;
wire
CORETSE_AHBiO10I
;
wire
CORETSE_AHBOI10I
;
assign
CORETSE_AHBoI1lI
=
CORETSE_AHBiII0I
;
assign
CORETSE_AHBiI1lI
=
CORETSE_AHBOIl0I
;
assign
CORETSE_AHBOl1lI
=
CORETSE_AHBlII0I
;
assign
CORETSE_AHBli1lI
=
CORETSE_AHBllI0I
;
assign
CORETSE_AHBll1lI
=
{
CORETSE_AHBO1olI
,
CORETSE_AHBo0olI
,
CORETSE_AHBI0olI
}
;
assign
CORETSE_AHBol1lI
=
{
CORETSE_AHBIoolI
,
CORETSE_AHBi1olI
,
CORETSE_AHBl1olI
}
;
assign
CORETSE_AHBil1lI
=
{
CORETSE_AHBliolI
,
CORETSE_AHBOiolI
,
CORETSE_AHBooolI
}
;
assign
CORETSE_AHBO01lI
=
CORETSE_AHBiiolI
;
assign
CORETSE_AHBI01lI
=
CORETSE_AHBIOilI
;
assign
CORETSE_AHBl01lI
=
CORETSE_AHBoOilI
;
assign
CORETSE_AHBOo1lI
=
CORETSE_AHBIol0I
;
assign
CORETSE_AHBo01lI
=
CORETSE_AHBolI0I
;
assign
CORETSE_AHBolI0I
=
CORETSE_AHBOIilI
[
`CORETSE_AHBoII0
]
;
assign
CORETSE_AHBi01lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBiII0
]
;
assign
CORETSE_AHBO11lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBOlI0
]
;
assign
CORETSE_AHBI11lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBIlI0
]
;
assign
CORETSE_AHBl11lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBllI0
]
;
assign
CORETSE_AHBo11lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBolI0
]
;
assign
CORETSE_AHBi11lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBilI0
]
;
assign
CORETSE_AHBio1lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBO0I0
]
;
assign
CORETSE_AHBOi1lI
=
CORETSE_AHBOIilI
[
`CORETSE_AHBI0I0
]
;
assign
CORETSE_AHBII10I
=
CORETSE_AHBOIilI
[
`CORETSE_AHBl0I0
]
;
assign
CORETSE_AHBlI10I
=
CORETSE_AHBOIilI
[
`CORETSE_AHBo0I0
]
;
assign
CORETSE_AHBoI10I
=
CORETSE_AHBOIilI
[
`CORETSE_AHBi0I0
]
;
assign
CORETSE_AHBlll0I
=
CORETSE_AHBOIilI
[
`CORETSE_AHBO1I0
]
;
assign
CORETSE_AHBIl1lI
=
CORETSE_AHBlll0I
;
assign
CORETSE_AHBIo1lI
=
CORETSE_AHBIlilI
;
assign
CORETSE_AHBlo1lI
=
CORETSE_AHBolilI
;
assign
CORETSE_AHBoo1lI
=
CORETSE_AHBOOI0I
;
assign
CORETSE_AHBIi1lI
=
CORETSE_AHBiOI0I
;
assign
CORETSE_AHBoi1lI
=
CORETSE_AHBO0I0I
;
assign
CORETSE_AHBii1lI
=
CORETSE_AHBloI0I
;
assign
CORETSE_AHBl0I0I
=
CORETSE_AHBO0I0I
&
~
CORETSE_AHBI0I0I
;
assign
CORETSE_AHBiI10I
=
CORETSE_AHBloI0I
&
~
CORETSE_AHBooI0I
;
assign
CORETSE_AHBOl10I
=
CORETSE_AHBlll0I
|
CORETSE_AHBi10lI
;
assign
CORETSE_AHBIoO0I
=
CORETSE_AHBIo0lI
;
assign
CORETSE_AHBIIl0I
=
~
CORETSE_AHBiIl0I
&
(
CORETSE_AHBIoO0I
|
(
~
CORETSE_AHBIoO0I
&
CORETSE_AHBlIl0I
)
)
;
assign
{
CORETSE_AHBO0olI
[
15
:
0
]
,
CORETSE_AHBololI
[
31
:
0
]
,
CORETSE_AHBIlolI
[
31
:
0
]
}
=
{
80
{
CORETSE_AHBIoO0I
}
}
&
CORETSE_AHBOi0lI
[
79
:
0
]
|
{
80
{
~
CORETSE_AHBIoO0I
}
}
&
{
CORETSE_AHBilolI
[
15
:
0
]
,
CORETSE_AHBllolI
[
31
:
0
]
,
CORETSE_AHBOlolI
[
31
:
0
]
}
;
assign
{
CORETSE_AHBiIolI
[
15
:
0
]
,
CORETSE_AHBlIolI
[
31
:
0
]
,
CORETSE_AHBOIolI
[
31
:
0
]
}
=
{
80
{
CORETSE_AHBOll0I
}
}
&
{
CORETSE_AHBilolI
[
15
:
0
]
,
CORETSE_AHBllolI
[
31
:
0
]
,
CORETSE_AHBOlolI
[
31
:
0
]
}
|
{
80
{
~
CORETSE_AHBOll0I
}
}
&
{
CORETSE_AHBoIolI
[
15
:
0
]
,
CORETSE_AHBIIolI
[
31
:
0
]
,
CORETSE_AHBiOolI
[
31
:
0
]
}
;
assign
CORETSE_AHBiOilI
=
(
CORETSE_AHBloO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBI1I0
]
|
~
(
CORETSE_AHBloO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBoOilI
&
~
CORETSE_AHBlOI0I
;
assign
CORETSE_AHBIIilI
=
{
(
`CORETSE_AHBO1I0
+
1
)
{
(
CORETSE_AHBooO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
`CORETSE_AHBO1I0
:
0
]
|
{
(
`CORETSE_AHBO1I0
+
1
)
{
~
(
CORETSE_AHBooO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBOIilI
;
assign
CORETSE_AHBoO10I
=
CORETSE_AHBOi00I
&
~
CORETSE_AHBIi00I
;
assign
CORETSE_AHBiO10I
=
CORETSE_AHBoi00I
&
~
CORETSE_AHBii00I
;
assign
CORETSE_AHBOI10I
=
CORETSE_AHBIO10I
&
~
CORETSE_AHBlO10I
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBl1O0
]
=
CORETSE_AHBOOI0I
|
~
CORETSE_AHBOOI0I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBl1O0
]
|
~
CORETSE_AHBOOI0I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBl1O0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBo1O0
]
=
CORETSE_AHBiOI0I
|
~
CORETSE_AHBiOI0I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBo1O0
]
|
~
CORETSE_AHBiOI0I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBo1O0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBi1O0
]
=
CORETSE_AHBlOI0I
|
~
CORETSE_AHBlOI0I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBi1O0
]
|
~
CORETSE_AHBlOI0I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBi1O0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBOoO0
]
=
CORETSE_AHBOOO0I
|
~
CORETSE_AHBOOO0I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBOoO0
]
|
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBOoO0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBIoO0
]
=
CORETSE_AHBI0O0I
|
~
CORETSE_AHBI0O0I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBIoO0
]
|
~
CORETSE_AHBI0O0I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBIoO0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBloO0
]
=
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBloO0
]
|
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBOII0I
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBooO0
]
=
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBooO0
]
|
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBIII0I
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBioO0
]
=
CORETSE_AHBoO10I
|
~
CORETSE_AHBoO10I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBioO0
]
|
~
CORETSE_AHBoO10I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBioO0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBOiO0
]
=
CORETSE_AHBiO10I
|
~
CORETSE_AHBiO10I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBOiO0
]
|
~
CORETSE_AHBiO10I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBOiO0
]
;
assign
CORETSE_AHBoIilI
[
`CORETSE_AHBIiO0
]
=
CORETSE_AHBOI10I
|
~
CORETSE_AHBOI10I
&
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBio0lI
[
`CORETSE_AHBIiO0
]
|
~
CORETSE_AHBOI10I
&
~
(
CORETSE_AHBOiO0I
&
~
CORETSE_AHBoo0lI
)
&
CORETSE_AHBlIilI
[
`CORETSE_AHBIiO0
]
;
assign
CORETSE_AHBOlilI
=
{
11
{
(
CORETSE_AHBioO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
10
:
0
]
|
{
11
{
~
(
CORETSE_AHBioO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBiIilI
;
assign
CORETSE_AHBl0olI
=
{
32
{
(
CORETSE_AHBIiO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
|
{
32
{
~
(
CORETSE_AHBIiO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBI0olI
;
assign
CORETSE_AHBi0olI
=
{
32
{
(
CORETSE_AHBliO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
|
{
32
{
~
(
CORETSE_AHBliO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBo0olI
;
assign
CORETSE_AHBI1olI
=
{
16
{
(
CORETSE_AHBoiO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
15
:
0
]
|
{
16
{
~
(
CORETSE_AHBoiO0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBO1olI
;
assign
CORETSE_AHBo1olI
=
{
32
{
(
CORETSE_AHBO0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
|
{
32
{
~
(
CORETSE_AHBO0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBl1olI
;
assign
CORETSE_AHBOoolI
=
{
32
{
(
CORETSE_AHBI0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
|
{
32
{
~
(
CORETSE_AHBI0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBi1olI
;
assign
CORETSE_AHBloolI
=
{
16
{
(
CORETSE_AHBl0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
15
:
0
]
|
{
16
{
~
(
CORETSE_AHBl0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBIoolI
;
assign
CORETSE_AHBOOilI
=
{
8
{
(
CORETSE_AHBo0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
7
:
0
]
|
{
8
{
~
(
CORETSE_AHBo0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBiiolI
;
assign
CORETSE_AHBioolI
=
{
32
{
(
CORETSE_AHBi0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
|
{
32
{
~
(
CORETSE_AHBi0ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBooolI
;
assign
CORETSE_AHBIiolI
=
{
32
{
(
CORETSE_AHBO1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
|
{
32
{
~
(
CORETSE_AHBO1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBOiolI
;
assign
CORETSE_AHBoiolI
=
{
16
{
(
CORETSE_AHBI1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
15
:
0
]
|
{
16
{
~
(
CORETSE_AHBI1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBliolI
;
assign
CORETSE_AHBlOilI
=
{
8
{
(
CORETSE_AHBl1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
7
:
0
]
|
{
8
{
~
(
CORETSE_AHBl1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBIOilI
;
assign
CORETSE_AHBllilI
=
{
(
CORETSE_AHBlII
-
CORETSE_AHBIII
+
1
)
{
(
CORETSE_AHBo1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
CORETSE_AHBlII
-
CORETSE_AHBIII
:
0
]
|
{
(
CORETSE_AHBlII
-
CORETSE_AHBIII
+
1
)
{
~
(
CORETSE_AHBo1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBIlilI
;
assign
CORETSE_AHBililI
=
{
(
CORETSE_AHBiII
-
CORETSE_AHBoII
+
1
)
{
(
CORETSE_AHBi1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
CORETSE_AHBiII
-
CORETSE_AHBoII
:
0
]
|
{
(
CORETSE_AHBiII
-
CORETSE_AHBoII
+
1
)
{
~
(
CORETSE_AHBi1ilI
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBolilI
;
assign
CORETSE_AHBlol0I
=
{
32
{
(
CORETSE_AHBi0l0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBio0lI
[
31
:
0
]
|
{
32
{
~
(
CORETSE_AHBi0l0I
&
~
CORETSE_AHBoo0lI
)
}
}
&
CORETSE_AHBIol0I
;
assign
CORETSE_AHBl000I
=
~
CORETSE_AHBi100I
&
(
CORETSE_AHBOI00I
|
CORETSE_AHBo000I
)
;
assign
CORETSE_AHBi000I
=
~
CORETSE_AHBIo00I
&
(
CORETSE_AHBII00I
|
CORETSE_AHBO100I
)
;
assign
CORETSE_AHBI100I
=
~
CORETSE_AHBoo00I
&
(
CORETSE_AHBlI00I
|
CORETSE_AHBl100I
)
;
assign
CORETSE_AHBOI00I
=
CORETSE_AHBiI00I
&
~
CORETSE_AHBOl00I
;
assign
CORETSE_AHBiol0I
=
{
32
{
(
CORETSE_AHBII10I
&
CORETSE_AHBOI00I
)
}
}
&
CORETSE_AHBOi0lI
[
31
:
0
]
|
{
32
{
~
(
CORETSE_AHBII10I
&
CORETSE_AHBOI00I
)
}
}
&
CORETSE_AHBool0I
;
assign
CORETSE_AHBIil0I
=
{
32
{
(
CORETSE_AHBII10I
&
CORETSE_AHBOI00I
)
}
}
&
CORETSE_AHBOi0lI
[
63
:
32
]
|
{
32
{
~
(
CORETSE_AHBII10I
&
CORETSE_AHBOI00I
)
}
}
&
CORETSE_AHBOil0I
;
assign
CORETSE_AHBII00I
=
CORETSE_AHBll00I
&
~
CORETSE_AHBol00I
;
assign
CORETSE_AHBoil0I
=
{
32
{
(
CORETSE_AHBlI10I
&
CORETSE_AHBII00I
)
}
}
&
CORETSE_AHBOi0lI
[
31
:
0
]
|
{
32
{
~
(
CORETSE_AHBlI10I
&
CORETSE_AHBII00I
)
}
}
&
CORETSE_AHBlil0I
;
assign
CORETSE_AHBOO00I
=
{
32
{
(
CORETSE_AHBlI10I
&
CORETSE_AHBII00I
)
}
}
&
CORETSE_AHBOi0lI
[
63
:
32
]
|
{
32
{
~
(
CORETSE_AHBlI10I
&
CORETSE_AHBII00I
)
}
}
&
CORETSE_AHBiil0I
;
assign
CORETSE_AHBlI00I
=
CORETSE_AHBO000I
&
~
CORETSE_AHBI000I
;
assign
CORETSE_AHBlO00I
=
{
32
{
(
CORETSE_AHBoI10I
&
CORETSE_AHBlI00I
)
}
}
&
CORETSE_AHBOi0lI
[
31
:
0
]
|
{
32
{
~
(
CORETSE_AHBoI10I
&
CORETSE_AHBlI00I
)
}
}
&
CORETSE_AHBIO00I
;
assign
CORETSE_AHBiO00I
=
{
32
{
(
CORETSE_AHBoI10I
&
CORETSE_AHBlI00I
)
}
}
&
CORETSE_AHBOi0lI
[
63
:
32
]
|
{
32
{
~
(
CORETSE_AHBoI10I
&
CORETSE_AHBlI00I
)
}
}
&
CORETSE_AHBoO00I
;
assign
CORETSE_AHBiII0I
[
31
:
0
]
=
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBlOl0I
)
}
}
&
CORETSE_AHBiOolI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBoOl0I
)
}
}
&
CORETSE_AHBIIolI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBiOl0I
)
}
}
&
{
16
'b
0
,
CORETSE_AHBoIolI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBloO0I
)
}
}
&
{
31
'b
0
,
CORETSE_AHBoOilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBooO0I
)
}
}
&
{
{
(
31
-
`CORETSE_AHBO1I0
)
{
1
'b
0
}
}
,
CORETSE_AHBOIilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBOiO0I
)
}
}
&
{
22
'b
0
,
CORETSE_AHBlIilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBioO0I
)
}
}
&
{
21
'b
0
,
CORETSE_AHBiIilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBIiO0I
)
}
}
&
CORETSE_AHBI0olI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBliO0I
)
}
}
&
CORETSE_AHBo0olI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBoiO0I
)
}
}
&
{
16
'b
0
,
CORETSE_AHBO1olI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBO0ilI
)
}
}
&
CORETSE_AHBl1olI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBI0ilI
)
}
}
&
CORETSE_AHBi1olI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBl0ilI
)
}
}
&
{
16
'b
0
,
CORETSE_AHBIoolI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBi0ilI
)
}
}
&
CORETSE_AHBooolI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBO1ilI
)
}
}
&
CORETSE_AHBOiolI
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBI1ilI
)
}
}
&
{
16
'b
0
,
CORETSE_AHBliolI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBo0ilI
)
}
}
&
{
24
'b
0
,
CORETSE_AHBiiolI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBl1ilI
)
}
}
&
{
24
'b
0
,
CORETSE_AHBIOilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBo1ilI
)
}
}
&
{
{
(
31
-
(
CORETSE_AHBlII
-
CORETSE_AHBIII
)
)
{
1
'b
0
}
}
,
CORETSE_AHBIlilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBi1ilI
)
}
}
&
{
{
(
31
-
(
CORETSE_AHBiII
-
CORETSE_AHBoII
)
)
{
1
'b
0
}
}
,
CORETSE_AHBolilI
}
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBIlI0I
)
}
}
&
CORETSE_AHBo1O0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBOlI0I
)
}
}
&
CORETSE_AHBOoO0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBi0l0I
)
}
}
&
CORETSE_AHBIol0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBO1l0I
)
}
}
&
CORETSE_AHBool0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBI1l0I
)
}
}
&
CORETSE_AHBOil0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBl1l0I
)
}
}
&
CORETSE_AHBlil0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBo1l0I
)
}
}
&
CORETSE_AHBiil0I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBi1l0I
)
}
}
&
CORETSE_AHBIO00I
|
{
32
{
(
CORETSE_AHBoo0lI
&
CORETSE_AHBOol0I
)
}
}
&
CORETSE_AHBoO00I
;
assign
CORETSE_AHBOIl0I
=
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBoII0I
=
CORETSE_AHBiIilI
[
`CORETSE_AHBliO0
]
&
(
(
CORETSE_AHBiIilI
[
`CORETSE_AHBoiO0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBl1O0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBiiO0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBo1O0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBOOI0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBi1O0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBIOI0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBOoO0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBlOI0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBIoO0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBoOI0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBloO0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBiOI0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBooO0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBOII0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBioO0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBIII0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBOiO0
]
)
|
(
CORETSE_AHBiIilI
[
`CORETSE_AHBlII0
]
&
CORETSE_AHBlIilI
[
`CORETSE_AHBIiO0
]
)
)
;
assign
CORETSE_AHBIoilI
=
(
~
CORETSE_AHBolI0I
|
(
~
CORETSE_AHBl0I0I
&
CORETSE_AHBOoilI
)
)
|
CORETSE_AHBOOO0I
;
assign
CORETSE_AHBooilI
=
CORETSE_AHBolI0I
&
CORETSE_AHBl0I0I
&
CORETSE_AHBOoilI
;
assign
CORETSE_AHBOiilI
=
CORETSE_AHBloilI
;
assign
CORETSE_AHBliilI
=
CORETSE_AHBioilI
;
assign
CORETSE_AHBiiilI
=
CORETSE_AHBIiilI
;
assign
CORETSE_AHBIOO0I
=
CORETSE_AHBoiilI
;
assign
CORETSE_AHBoOO0I
=
(
CORETSE_AHBolI0I
&
CORETSE_AHBl0I0I
&
CORETSE_AHBOoilI
)
|
CORETSE_AHBloilI
|
CORETSE_AHBioilI
|
CORETSE_AHBIiilI
|
CORETSE_AHBoiilI
|
CORETSE_AHBOOO0I
;
assign
CORETSE_AHBOIO0I
[
0
]
=
CORETSE_AHBolI0I
&
CORETSE_AHBl0I0I
&
CORETSE_AHBOoilI
;
assign
CORETSE_AHBOIO0I
[
1
]
=
CORETSE_AHBloilI
;
assign
CORETSE_AHBOIO0I
[
2
]
=
CORETSE_AHBioilI
;
assign
CORETSE_AHBOIO0I
[
3
]
=
CORETSE_AHBIiilI
;
assign
CORETSE_AHBOIO0I
[
4
]
=
CORETSE_AHBoiilI
;
assign
CORETSE_AHBOIO0I
[
5
]
=
CORETSE_AHBOOO0I
;
assign
CORETSE_AHBl1O0I
=
(
{
32
{
CORETSE_AHBiOO0I
[
0
]
}
}
&
{
CORETSE_AHBo0I0I
[
15
:
0
]
,
12
'b
0
,
CORETSE_AHBO1I0I
[
3
:
0
]
}
)
|
(
{
32
{
CORETSE_AHBiOO0I
[
1
]
}
}
&
CORETSE_AHBl1I0I
[
31
:
0
]
)
|
(
{
32
{
CORETSE_AHBiOO0I
[
2
]
}
}
&
CORETSE_AHBl1I0I
[
63
:
32
]
)
|
(
{
32
{
CORETSE_AHBiOO0I
[
3
]
}
}
&
{
CORETSE_AHBi1I0I
[
15
:
0
]
,
CORETSE_AHBl1I0I
[
79
:
64
]
}
)
|
(
{
32
{
CORETSE_AHBiOO0I
[
4
]
}
}
&
CORETSE_AHBi1I0I
[
47
:
16
]
)
|
(
{
32
{
CORETSE_AHBiOO0I
[
5
]
}
}
&
CORETSE_AHBi1I0I
[
79
:
48
]
)
;
assign
CORETSE_AHBi0I0I
=
{
16
{
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBlO1lI
|
{
16
{
~
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBo0I0I
;
assign
CORETSE_AHBI1I0I
=
{
4
{
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBIO1lI
|
{
4
{
~
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBO1I0I
;
assign
CORETSE_AHBo1I0I
=
{
80
{
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBoO1lI
|
{
80
{
~
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBl1I0I
;
assign
CORETSE_AHBOoI0I
=
{
80
{
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBioo1
|
{
80
{
~
CORETSE_AHBl0I0I
}
}
&
CORETSE_AHBi1I0I
;
assign
CORETSE_AHBlIO0I
=
(
~
CORETSE_AHBolI0I
|
(
~
CORETSE_AHBiI10I
&
CORETSE_AHBIIO0I
)
)
|
CORETSE_AHBI0O0I
;
assign
CORETSE_AHBiIO0I
=
CORETSE_AHBolI0I
&
CORETSE_AHBiI10I
&
CORETSE_AHBIIO0I
;
assign
CORETSE_AHBIlO0I
=
CORETSE_AHBoIO0I
;
assign
CORETSE_AHBolO0I
=
CORETSE_AHBOlO0I
;
assign
CORETSE_AHBO0O0I
=
CORETSE_AHBllO0I
;
assign
CORETSE_AHBl0O0I
=
CORETSE_AHBilO0I
;
assign
CORETSE_AHBi0O0I
=
(
CORETSE_AHBolI0I
&
CORETSE_AHBiI10I
&
CORETSE_AHBIIO0I
)
|
CORETSE_AHBoIO0I
|
CORETSE_AHBOlO0I
|
CORETSE_AHBllO0I
|
CORETSE_AHBilO0I
|
CORETSE_AHBI0O0I
;
assign
CORETSE_AHBI1O0I
[
0
]
=
CORETSE_AHBolI0I
&
CORETSE_AHBiI10I
&
CORETSE_AHBIIO0I
;
assign
CORETSE_AHBI1O0I
[
1
]
=
CORETSE_AHBoIO0I
;
assign
CORETSE_AHBI1O0I
[
2
]
=
CORETSE_AHBOlO0I
;
assign
CORETSE_AHBI1O0I
[
3
]
=
CORETSE_AHBllO0I
;
assign
CORETSE_AHBI1O0I
[
4
]
=
CORETSE_AHBilO0I
;
assign
CORETSE_AHBI1O0I
[
5
]
=
CORETSE_AHBI0O0I
;
assign
CORETSE_AHBi1O0I
=
{
32
{
CORETSE_AHBO1O0I
[
0
]
}
}
&
(
{
CORETSE_AHBioI0I
[
15
:
0
]
,
12
'b
000000000000
,
CORETSE_AHBIiI0I
[
3
:
0
]
}
)
|
{
32
{
CORETSE_AHBO1O0I
[
1
]
}
}
&
CORETSE_AHBoiI0I
[
31
:
0
]
|
{
32
{
CORETSE_AHBO1O0I
[
2
]
}
}
&
CORETSE_AHBoiI0I
[
63
:
32
]
|
{
32
{
CORETSE_AHBO1O0I
[
3
]
}
}
&
(
{
CORETSE_AHBOOl0I
[
15
:
0
]
,
CORETSE_AHBoiI0I
[
79
:
64
]
}
)
|
{
32
{
CORETSE_AHBO1O0I
[
4
]
}
}
&
CORETSE_AHBOOl0I
[
47
:
16
]
|
{
32
{
CORETSE_AHBO1O0I
[
5
]
}
}
&
CORETSE_AHBOOl0I
[
79
:
48
]
;
assign
CORETSE_AHBOiI0I
=
{
16
{
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBOI1lI
|
{
16
{
~
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBioI0I
;
assign
CORETSE_AHBliI0I
=
{
4
{
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBiO1lI
|
{
4
{
~
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBIiI0I
;
assign
CORETSE_AHBiiI0I
=
{
80
{
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBII1lI
|
{
80
{
~
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBoiI0I
;
assign
CORETSE_AHBIOl0I
=
{
80
{
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBlI1lI
|
{
80
{
~
CORETSE_AHBiI10I
}
}
&
CORETSE_AHBOOl0I
;
assign
CORETSE_AHBO0l0I
=
CORETSE_AHBill0I
&
CORETSE_AHBlOO0I
&
~
CORETSE_AHBl0l0I
;
assign
CORETSE_AHBI0l0I
=
CORETSE_AHBoll0I
&
CORETSE_AHBo0O0I
&
~
CORETSE_AHBo0l0I
;
sib_fifo_top
#
(
.CORETSE_AHBIl10I
(
32
)
,
.CORETSE_AHBll10I
(
CORETSE_AHBllI
)
,
.CORETSE_AHBol10I
(
0
)
,
.CORETSE_AHBil10I
(
0
)
,
.CORETSE_AHBO010I
(
0
)
,
.CORETSE_AHBI010I
(
0
)
)
CORETSE_AHBl010I
(
.CORETSE_AHBo010I
(
CORETSE_AHBiil0
)
,
.CORETSE_AHBi010I
(
~
CORETSE_AHBOl10I
)
,
.CORETSE_AHBO110I
(
CORETSE_AHBiil0
)
,
.CORETSE_AHBI110I
(
~
CORETSE_AHBOl10I
)
,
.CORETSE_AHBl110I
(
CORETSE_AHBl1O0I
)
,
.CORETSE_AHBo110I
(
CORETSE_AHBo1O0I
)
,
.CORETSE_AHBi110I
(
CORETSE_AHBO0l0I
)
,
.CORETSE_AHBOo10I
(
CORETSE_AHBOOolI
)
,
.CORETSE_AHBIo10I
(
CORETSE_AHBl0l0I
)
,
.CORETSE_AHBlo10I
(
CORETSE_AHBOII0I
)
,
.CORETSE_AHBoo10I
(
)
,
.CORETSE_AHBio10I
(
)
,
.CORETSE_AHBOi10I
(
CORETSE_AHBIlI0I
&
CORETSE_AHBoo0lI
)
,
.CORETSE_AHBIi10I
(
CORETSE_AHBlOolI
)
,
.CORETSE_AHBli10I
(
)
,
.CORETSE_AHBoi10I
(
CORETSE_AHBill0I
)
)
;
sib_fifo_top
#
(
.CORETSE_AHBIl10I
(
32
)
,
.CORETSE_AHBll10I
(
CORETSE_AHBolI
)
,
.CORETSE_AHBol10I
(
0
)
,
.CORETSE_AHBil10I
(
0
)
,
.CORETSE_AHBO010I
(
0
)
,
.CORETSE_AHBI010I
(
0
)
)
CORETSE_AHBii10I
(
.CORETSE_AHBo010I
(
CORETSE_AHBiil0
)
,
.CORETSE_AHBi010I
(
~
CORETSE_AHBOl10I
)
,
.CORETSE_AHBO110I
(
CORETSE_AHBiil0
)
,
.CORETSE_AHBI110I
(
~
CORETSE_AHBOl10I
)
,
.CORETSE_AHBl110I
(
CORETSE_AHBi1O0I
)
,
.CORETSE_AHBo110I
(
CORETSE_AHBOoO0I
)
,
.CORETSE_AHBi110I
(
CORETSE_AHBI0l0I
)
,
.CORETSE_AHBOo10I
(
CORETSE_AHBIOolI
)
,
.CORETSE_AHBIo10I
(
CORETSE_AHBo0l0I
)
,
.CORETSE_AHBlo10I
(
CORETSE_AHBIII0I
)
,
.CORETSE_AHBoo10I
(
)
,
.CORETSE_AHBio10I
(
)
,
.CORETSE_AHBOi10I
(
CORETSE_AHBOlI0I
&
CORETSE_AHBoo0lI
)
,
.CORETSE_AHBIi10I
(
CORETSE_AHBoOolI
)
,
.CORETSE_AHBli10I
(
)
,
.CORETSE_AHBoi10I
(
CORETSE_AHBoll0I
)
)
;
assign
CORETSE_AHBlOl0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBooil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBoOl0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBioil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBiOl0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBOiil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBIiO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBIiil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBliO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBliil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBoiO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBoiil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBO0ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBiiil
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBI0ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBOOO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBl0ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBIOO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBi0ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBlOO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBO1ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBoOO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBI1ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBiOO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBo0ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBOIO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBl1ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBIIO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBloO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBlIO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBooO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBoIO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBOiO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBiIO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBioO0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBOlO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBo1ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBIlO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBi1ilI
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBllO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBOlI0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBolO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBIlI0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBilO0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBi0l0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBO0O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBO1l0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBI0O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBI1l0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBl0O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBl1l0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBo0O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBo1l0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBi0O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBi1l0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBO1O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBOol0I
=
(
CORETSE_AHBoO00
==
`CORETSE_AHBI1O0
)
&
~
CORETSE_AHBlo0lI
;
assign
CORETSE_AHBllI0I
=
~
CORETSE_AHBlo0lI
&
CORETSE_AHBoo0lI
;
always
@
(
posedge
CORETSE_AHBiil0
or
posedge
CORETSE_AHBi10lI
)
begin
if
(
CORETSE_AHBi10lI
)
begin
CORETSE_AHBI0olI
<=
32
'b
0
;
CORETSE_AHBo0olI
<=
32
'b
0
;
CORETSE_AHBO1olI
<=
16
'b
0
;
CORETSE_AHBoOilI
<=
1
'b
0
;
CORETSE_AHBOIilI
<=
{
(
`CORETSE_AHBO1I0
+
1
)
{
1
'b
0
}
}
;
CORETSE_AHBlIilI
<=
10
'b
0
;
CORETSE_AHBiIilI
<=
11
'b
0
;
CORETSE_AHBlII0I
<=
1
'b
0
;
CORETSE_AHBl1olI
<=
32
'b
0
;
CORETSE_AHBi1olI
<=
32
'b
0
;
CORETSE_AHBIoolI
<=
16
'b
0
;
CORETSE_AHBiiolI
<=
8
'b
00000001
;
CORETSE_AHBooolI
<=
32
'b
0
;
CORETSE_AHBOiolI
<=
32
'b
0
;
CORETSE_AHBliolI
<=
16
'b
0
;
CORETSE_AHBIOilI
<=
8
'b
00000001
;
CORETSE_AHBIlilI
<=
{
(
CORETSE_AHBlII
-
CORETSE_AHBIII
+
1
)
{
1
'b
0
}
}
;
CORETSE_AHBolilI
<=
{
(
CORETSE_AHBiII
-
CORETSE_AHBoII
+
1
)
{
1
'b
0
}
}
;
CORETSE_AHBiOolI
<=
32
'b
0
;
CORETSE_AHBIIolI
<=
32
'b
0
;
CORETSE_AHBoIolI
<=
16
'b
0
;
CORETSE_AHBIol0I
<=
32
'b
0
;
end
else
begin
CORETSE_AHBI0olI
<=
CORETSE_AHBl0olI
;
CORETSE_AHBo0olI
<=
CORETSE_AHBi0olI
;
CORETSE_AHBO1olI
<=
CORETSE_AHBI1olI
;
CORETSE_AHBoOilI
<=
CORETSE_AHBiOilI
;
CORETSE_AHBOIilI
<=
CORETSE_AHBIIilI
;
CORETSE_AHBlIilI
<=
CORETSE_AHBoIilI
;
CORETSE_AHBiIilI
<=
CORETSE_AHBOlilI
;
CORETSE_AHBlII0I
<=
CORETSE_AHBoII0I
;
CORETSE_AHBl1olI
<=
CORETSE_AHBo1olI
;
CORETSE_AHBi1olI
<=
CORETSE_AHBOoolI
;
CORETSE_AHBIoolI
<=
CORETSE_AHBloolI
;
CORETSE_AHBiiolI
<=
CORETSE_AHBOOilI
;
CORETSE_AHBooolI
<=
CORETSE_AHBioolI
;
CORETSE_AHBOiolI
<=
CORETSE_AHBIiolI
;
CORETSE_AHBliolI
<=
CORETSE_AHBoiolI
;
CORETSE_AHBIOilI
<=
CORETSE_AHBlOilI
;
CORETSE_AHBIlilI
<=
CORETSE_AHBllilI
;
CORETSE_AHBolilI
<=
CORETSE_AHBililI
;
CORETSE_AHBiOolI
<=
CORETSE_AHBOIolI
;
CORETSE_AHBIIolI
<=
CORETSE_AHBlIolI
;
CORETSE_AHBoIolI
<=
CORETSE_AHBiIolI
;
CORETSE_AHBIol0I
<=
CORETSE_AHBlol0I
;
end
end
always
@
(
posedge
CORETSE_AHBiil0
or
posedge
CORETSE_AHBOl10I
)
begin
if
(
CORETSE_AHBOl10I
)
begin
CORETSE_AHBiiO0I
<=
1
'b
0
;
CORETSE_AHBOOI0I
<=
1
'b
0
;
CORETSE_AHBIOI0I
<=
1
'b
0
;
CORETSE_AHBlOI0I
<=
1
'b
0
;
CORETSE_AHBoOI0I
<=
1
'b
0
;
CORETSE_AHBiOI0I
<=
1
'b
0
;
CORETSE_AHBilI0I
<=
1
'b
0
;
CORETSE_AHBO0I0I
<=
1
'b
0
;
CORETSE_AHBI0I0I
<=
1
'b
0
;
CORETSE_AHBo0I0I
<=
16
'b
0
;
CORETSE_AHBO1I0I
<=
4
'b
0
;
CORETSE_AHBl1I0I
<=
80
'b
0
;
CORETSE_AHBi1I0I
<=
80
'b
0
;
CORETSE_AHBIoI0I
<=
1
'b
0
;
CORETSE_AHBloI0I
<=
1
'b
0
;
CORETSE_AHBooI0I
<=
1
'b
0
;
CORETSE_AHBioI0I
<=
16
'b
0
;
CORETSE_AHBIiI0I
<=
4
'b
0
;
CORETSE_AHBoiI0I
<=
80
'b
0
;
CORETSE_AHBOOl0I
<=
80
'b
0
;
CORETSE_AHBOoilI
<=
1
'b
0
;
CORETSE_AHBloilI
<=
1
'b
0
;
CORETSE_AHBioilI
<=
1
'b
0
;
CORETSE_AHBIiilI
<=
1
'b
0
;
CORETSE_AHBoiilI
<=
1
'b
0
;
CORETSE_AHBOOO0I
<=
1
'b
0
;
CORETSE_AHBlOO0I
<=
1
'b
0
;
CORETSE_AHBiOO0I
<=
6
'b
0
;
CORETSE_AHBIIO0I
<=
1
'b
0
;
CORETSE_AHBoIO0I
<=
1
'b
0
;
CORETSE_AHBOlO0I
<=
1
'b
0
;
CORETSE_AHBllO0I
<=
1
'b
0
;
CORETSE_AHBilO0I
<=
1
'b
0
;
CORETSE_AHBI0O0I
<=
1
'b
0
;
CORETSE_AHBo0O0I
<=
1
'b
0
;
CORETSE_AHBO1O0I
<=
6
'b
0
;
CORETSE_AHBIll0I
<=
1
'b
0
;
CORETSE_AHBOll0I
<=
1
'b
0
;
CORETSE_AHBio00I
<=
1
'b
0
;
CORETSE_AHBOi00I
<=
1
'b
0
;
CORETSE_AHBIi00I
<=
1
'b
0
;
CORETSE_AHBli00I
<=
1
'b
0
;
CORETSE_AHBoi00I
<=
1
'b
0
;
CORETSE_AHBii00I
<=
1
'b
0
;
CORETSE_AHBOO10I
<=
1
'b
0
;
CORETSE_AHBIO10I
<=
1
'b
0
;
CORETSE_AHBlO10I
<=
1
'b
0
;
end
else
begin
CORETSE_AHBiiO0I
<=
CORETSE_AHBIi0lI
;
CORETSE_AHBOOI0I
<=
CORETSE_AHBiiO0I
;
CORETSE_AHBIOI0I
<=
CORETSE_AHBoi0lI
;
CORETSE_AHBlOI0I
<=
CORETSE_AHBIOI0I
;
CORETSE_AHBoOI0I
<=
CORETSE_AHBli0lI
;
CORETSE_AHBiOI0I
<=
CORETSE_AHBoOI0I
;
CORETSE_AHBilI0I
<=
CORETSE_AHBii0lI
;
CORETSE_AHBO0I0I
<=
CORETSE_AHBilI0I
;
CORETSE_AHBI0I0I
<=
CORETSE_AHBO0I0I
;
CORETSE_AHBo0I0I
<=
CORETSE_AHBi0I0I
;
CORETSE_AHBO1I0I
<=
CORETSE_AHBI1I0I
;
CORETSE_AHBl1I0I
<=
CORETSE_AHBo1I0I
;
CORETSE_AHBi1I0I
<=
CORETSE_AHBOoI0I
;
CORETSE_AHBIoI0I
<=
CORETSE_AHBOO1lI
;
CORETSE_AHBloI0I
<=
CORETSE_AHBIoI0I
;
CORETSE_AHBooI0I
<=
CORETSE_AHBloI0I
;
CORETSE_AHBioI0I
<=
CORETSE_AHBOiI0I
;
CORETSE_AHBIiI0I
<=
CORETSE_AHBliI0I
;
CORETSE_AHBoiI0I
<=
CORETSE_AHBiiI0I
;
CORETSE_AHBOOl0I
<=
CORETSE_AHBIOl0I
;
CORETSE_AHBOoilI
<=
CORETSE_AHBIoilI
;
CORETSE_AHBloilI
<=
CORETSE_AHBooilI
;
CORETSE_AHBioilI
<=
CORETSE_AHBOiilI
;
CORETSE_AHBIiilI
<=
CORETSE_AHBliilI
;
CORETSE_AHBoiilI
<=
CORETSE_AHBiiilI
;
CORETSE_AHBOOO0I
<=
CORETSE_AHBIOO0I
;
CORETSE_AHBlOO0I
<=
CORETSE_AHBoOO0I
;
CORETSE_AHBiOO0I
<=
CORETSE_AHBOIO0I
;
CORETSE_AHBIIO0I
<=
CORETSE_AHBlIO0I
;
CORETSE_AHBoIO0I
<=
CORETSE_AHBiIO0I
;
CORETSE_AHBOlO0I
<=
CORETSE_AHBIlO0I
;
CORETSE_AHBllO0I
<=
CORETSE_AHBolO0I
;
CORETSE_AHBilO0I
<=
CORETSE_AHBO0O0I
;
CORETSE_AHBI0O0I
<=
CORETSE_AHBl0O0I
;
CORETSE_AHBo0O0I
<=
CORETSE_AHBi0O0I
;
CORETSE_AHBO1O0I
<=
CORETSE_AHBI1O0I
;
CORETSE_AHBIll0I
<=
CORETSE_AHBlIl0I
;
CORETSE_AHBOll0I
<=
CORETSE_AHBIll0I
;
CORETSE_AHBio00I
<=
CORETSE_AHBo000I
;
CORETSE_AHBOi00I
<=
CORETSE_AHBio00I
;
CORETSE_AHBIi00I
<=
CORETSE_AHBOi00I
;
CORETSE_AHBli00I
<=
CORETSE_AHBO100I
;
CORETSE_AHBoi00I
<=
CORETSE_AHBli00I
;
CORETSE_AHBii00I
<=
CORETSE_AHBoi00I
;
CORETSE_AHBOO10I
<=
CORETSE_AHBl100I
;
CORETSE_AHBIO10I
<=
CORETSE_AHBOO10I
;
CORETSE_AHBlO10I
<=
CORETSE_AHBIO10I
;
end
end
always
@
(
posedge
CORETSE_AHBOl0
or
posedge
CORETSE_AHBOo0lI
)
begin
if
(
CORETSE_AHBOo0lI
)
begin
CORETSE_AHBoIl0I
<=
1
'b
0
;
CORETSE_AHBiIl0I
<=
1
'b
0
;
CORETSE_AHBOlolI
<=
32
'b
0
;
CORETSE_AHBllolI
<=
32
'b
0
;
CORETSE_AHBilolI
<=
16
'b
0
;
CORETSE_AHBlIl0I
<=
1
'b
0
;
CORETSE_AHBool0I
<=
32
'b
0
;
CORETSE_AHBOil0I
<=
32
'b
0
;
CORETSE_AHBlil0I
<=
32
'b
0
;
CORETSE_AHBiil0I
<=
32
'b
0
;
CORETSE_AHBIO00I
<=
32
'b
0
;
CORETSE_AHBoO00I
<=
32
'b
0
;
CORETSE_AHBoI00I
<=
1
'b
0
;
CORETSE_AHBiI00I
<=
1
'b
0
;
CORETSE_AHBOl00I
<=
1
'b
0
;
CORETSE_AHBIl00I
<=
1
'b
0
;
CORETSE_AHBll00I
<=
1
'b
0
;
CORETSE_AHBol00I
<=
1
'b
0
;
CORETSE_AHBil00I
<=
1
'b
0
;
CORETSE_AHBO000I
<=
1
'b
0
;
CORETSE_AHBI000I
<=
1
'b
0
;
CORETSE_AHBo000I
<=
1
'b
0
;
CORETSE_AHBO100I
<=
1
'b
0
;
CORETSE_AHBl100I
<=
1
'b
0
;
CORETSE_AHBo100I
<=
1
'b
0
;
CORETSE_AHBi100I
<=
1
'b
0
;
CORETSE_AHBOo00I
<=
1
'b
0
;
CORETSE_AHBIo00I
<=
1
'b
0
;
CORETSE_AHBlo00I
<=
1
'b
0
;
CORETSE_AHBoo00I
<=
1
'b
0
;
end
else
begin
CORETSE_AHBoIl0I
<=
CORETSE_AHBOll0I
;
CORETSE_AHBiIl0I
<=
CORETSE_AHBoIl0I
;
CORETSE_AHBOlolI
<=
CORETSE_AHBIlolI
;
CORETSE_AHBllolI
<=
CORETSE_AHBololI
;
CORETSE_AHBilolI
<=
CORETSE_AHBO0olI
;
CORETSE_AHBlIl0I
<=
CORETSE_AHBIIl0I
;
CORETSE_AHBool0I
<=
CORETSE_AHBiol0I
;
CORETSE_AHBOil0I
<=
CORETSE_AHBIil0I
;
CORETSE_AHBlil0I
<=
CORETSE_AHBoil0I
;
CORETSE_AHBiil0I
<=
CORETSE_AHBOO00I
;
CORETSE_AHBIO00I
<=
CORETSE_AHBlO00I
;
CORETSE_AHBoO00I
<=
CORETSE_AHBiO00I
;
CORETSE_AHBoI00I
<=
CORETSE_AHBlI0
;
CORETSE_AHBiI00I
<=
CORETSE_AHBoI00I
;
CORETSE_AHBOl00I
<=
CORETSE_AHBiI00I
;
CORETSE_AHBIl00I
<=
CORETSE_AHBoI0
;
CORETSE_AHBll00I
<=
CORETSE_AHBIl00I
;
CORETSE_AHBol00I
<=
CORETSE_AHBll00I
;
CORETSE_AHBil00I
<=
CORETSE_AHBiI0
;
CORETSE_AHBO000I
<=
CORETSE_AHBil00I
;
CORETSE_AHBI000I
<=
CORETSE_AHBO000I
;
CORETSE_AHBo000I
<=
CORETSE_AHBl000I
;
CORETSE_AHBO100I
<=
CORETSE_AHBi000I
;
CORETSE_AHBl100I
<=
CORETSE_AHBI100I
;
CORETSE_AHBo100I
<=
CORETSE_AHBOi00I
;
CORETSE_AHBi100I
<=
CORETSE_AHBo100I
;
CORETSE_AHBOo00I
<=
CORETSE_AHBoi00I
;
CORETSE_AHBIo00I
<=
CORETSE_AHBOo00I
;
CORETSE_AHBlo00I
<=
CORETSE_AHBIO10I
;
CORETSE_AHBoo00I
<=
CORETSE_AHBlo00I
;
end
end
endmodule
