//                        Proprietary and Confidential                          
//                  Copyright (c) 2013 All Rights Reserved                     
// REVISION    : $Revision: 1.5 $                                                  
module
sib_sync_2flp
#
(
parameter
CORETSE_AHBlIloI
=
1
,
parameter
CORETSE_AHBoIloI
=
0
)
(
input
CORETSE_AHBOlloI,
input
CORETSE_AHBIlloI,
input
CORETSE_AHBllloI,
input
CORETSE_AHBolloI,
input
[
CORETSE_AHBlIloI
-
1
:
0
]
CORETSE_AHBilloI,
output
[
CORETSE_AHBlIloI
-
1
:
0
]
CORETSE_AHBO0loI
)
;
reg
[
CORETSE_AHBlIloI
-
1
:
0
]
CORETSE_AHBl1loI
,
CORETSE_AHBo1loI
,
CORETSE_AHBi1loI
;
integer
CORETSE_AHBOloI
;
generate
if
(
CORETSE_AHBoIloI
==
1
)
begin
:
CORETSE_AHBOoloI
always
@
(
posedge
CORETSE_AHBOlloI
or
negedge
CORETSE_AHBllloI
)
begin
if
(
~
CORETSE_AHBllloI
)
CORETSE_AHBi1loI
<=
0
;
else
CORETSE_AHBi1loI
<=
CORETSE_AHBilloI
;
end
always
@
(
posedge
CORETSE_AHBIlloI
or
negedge
CORETSE_AHBolloI
)
begin
if
(
~
CORETSE_AHBolloI
)
begin
CORETSE_AHBl1loI
<=
0
;
CORETSE_AHBo1loI
<=
0
;
end
else
begin
CORETSE_AHBl1loI
<=
CORETSE_AHBi1loI
;
CORETSE_AHBo1loI
<=
CORETSE_AHBl1loI
;
end
end
end
else
begin
:
CORETSE_AHBIoloI
always
@
(
posedge
CORETSE_AHBOlloI
)
CORETSE_AHBi1loI
<=
CORETSE_AHBilloI
;
always
@
(
posedge
CORETSE_AHBIlloI
)
begin
CORETSE_AHBl1loI
<=
CORETSE_AHBi1loI
;
CORETSE_AHBo1loI
<=
CORETSE_AHBl1loI
;
end
end
endgenerate
assign
CORETSE_AHBO0loI
=
CORETSE_AHBo1loI
;
endmodule
