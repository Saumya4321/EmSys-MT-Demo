//                        Proprietary and Confidential                          
//                  Copyright (c) 2013 All Rights Reserved                     
// REVISION    : $Revision: 1.2 $                                                  
module
sib_fifo_mem2p
#
(
parameter
CORETSE_AHBIl10I
=
64
,
parameter
CORETSE_AHBol10I
=
0
,
parameter
CORETSE_AHBil10I
=
0
,
parameter
CORETSE_AHBO010I
=
0
,
parameter
CORETSE_AHBll10I
=
4
)
(
input
CORETSE_AHBo010I,
input
CORETSE_AHBO110I,
input
CORETSE_AHBI0IoI,
input
CORETSE_AHBl0IoI,
input
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBo0IoI,
input
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBi0IoI,
input
[
CORETSE_AHBIl10I
-
1
:
0
]
CORETSE_AHBl110I,
output
[
CORETSE_AHBIl10I
-
1
:
0
]
CORETSE_AHBo110I
)
;
localparam
CORETSE_AHBO1IoI
=
(
1
<<
CORETSE_AHBll10I
)
;
reg
[
CORETSE_AHBIl10I
-
1
:
0
]
CORETSE_AHBI1IoI
[
0
:
CORETSE_AHBO1IoI
-
1
]
;
reg
[
CORETSE_AHBll10I
-
1
:
0
]
CORETSE_AHBl1IoI
;
generate
integer
CORETSE_AHBOloI
;
if
(
CORETSE_AHBO010I
==
1
)
initial
for
(
CORETSE_AHBOloI
=
0
;
CORETSE_AHBOloI
<
CORETSE_AHBO1IoI
;
CORETSE_AHBOloI
=
CORETSE_AHBOloI
+
1
)
CORETSE_AHBI1IoI
[
CORETSE_AHBOloI
]
=
{
CORETSE_AHBIl10I
{
1
'b
0
}
}
;
endgenerate
assign
CORETSE_AHBo110I
=
CORETSE_AHBI1IoI
[
CORETSE_AHBl1IoI
]
;
generate
if
(
CORETSE_AHBil10I
==
1
)
always
@
(
posedge
CORETSE_AHBO110I
)
CORETSE_AHBl1IoI
<=
CORETSE_AHBl0IoI
?
CORETSE_AHBi0IoI
:
CORETSE_AHBl1IoI
;
else
if
(
CORETSE_AHBol10I
==
1
)
always
@
(
posedge
CORETSE_AHBO110I
)
CORETSE_AHBl1IoI
<=
CORETSE_AHBi0IoI
;
else
always
@
(
*
)
CORETSE_AHBl1IoI
=
CORETSE_AHBi0IoI
;
endgenerate
always
@
(
posedge
CORETSE_AHBo010I
)
begin
CORETSE_AHBI1IoI
[
CORETSE_AHBo0IoI
]
<=
CORETSE_AHBI0IoI
?
CORETSE_AHBl110I
:
CORETSE_AHBI1IoI
[
CORETSE_AHBo0IoI
]
;
end
endmodule
