`timescale 1 ns/100 ps
// Version: v11.7 SP2 11.7.2.2


module CoreTSE_Webserver_FCCC_3_FCCC(
       NGMUX0_SEL,
       NGMUX0_ARST_N,
       NGMUX0_HOLD_N,
       NGMUX1_SEL,
       NGMUX1_ARST_N,
       NGMUX1_HOLD_N,
       LOCK,
       CLK0,
       CLK1,
       GL0,
       GL1
    );
input  NGMUX0_SEL;
input  NGMUX0_ARST_N;
input  NGMUX0_HOLD_N;
input  NGMUX1_SEL;
input  NGMUX1_ARST_N;
input  NGMUX1_HOLD_N;
output LOCK;
input  CLK0;
input  CLK1;
output GL0;
output GL1;

    wire gnd_net, vcc_net, GL0_net, GL1_net;
    
    CLKINT GL1_INST (.A(GL1_net), .Y(GL1));
    VCC vcc_inst (.Y(vcc_net));
    GND gnd_inst (.Y(gnd_net));
    CLKINT GL0_INST (.A(GL0_net), .Y(GL0));
    CCC #( .INIT(210'h000C007FC0000044964001F18C613542B0739DF00404C81400303)
        , .VCOFREQUENCY(500.000) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(
        ), .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(
        LOCK), .BUSY(), .CLK0(CLK0), .CLK1(CLK1), .CLK2(vcc_net), 
        .CLK3(vcc_net), .NGMUX0_SEL(NGMUX0_SEL), .NGMUX1_SEL(
        NGMUX1_SEL), .NGMUX2_SEL(gnd_net), .NGMUX3_SEL(gnd_net), 
        .NGMUX0_HOLD_N(NGMUX0_HOLD_N), .NGMUX1_HOLD_N(NGMUX1_HOLD_N), 
        .NGMUX2_HOLD_N(vcc_net), .NGMUX3_HOLD_N(vcc_net), 
        .NGMUX0_ARST_N(NGMUX0_ARST_N), .NGMUX1_ARST_N(NGMUX1_ARST_N), 
        .NGMUX2_ARST_N(vcc_net), .NGMUX3_ARST_N(vcc_net), 
        .PLL_BYPASS_N(vcc_net), .PLL_ARST_N(vcc_net), .PLL_POWERDOWN_N(
        vcc_net), .GPD0_ARST_N(vcc_net), .GPD1_ARST_N(vcc_net), 
        .GPD2_ARST_N(vcc_net), .GPD3_ARST_N(vcc_net), .PRESET_N(
        gnd_net), .PCLK(vcc_net), .PSEL(vcc_net), .PENABLE(vcc_net), 
        .PWRITE(vcc_net), .PADDR({vcc_net, vcc_net, vcc_net, vcc_net, 
        vcc_net, vcc_net}), .PWDATA({vcc_net, vcc_net, vcc_net, 
        vcc_net, vcc_net, vcc_net, vcc_net, vcc_net}), .CLK0_PAD(
        gnd_net), .CLK1_PAD(gnd_net), .CLK2_PAD(gnd_net), .CLK3_PAD(
        gnd_net), .GL0(GL0_net), .GL1(GL1_net), .GL2(), .GL3(), 
        .RCOSC_25_50MHZ(gnd_net), .RCOSC_1MHZ(gnd_net), .XTLOSC(
        gnd_net));
    
endmodule
