//                        Proprietary and Confidential 
// REVISION    : $Revision: $ 
`include "include.v"
module
ptp_rfp
(
input
CORETSE_AHBOOo0I,
input
CORETSE_AHBIOo0I,
input
CORETSE_AHBlOo0I,
input
CORETSE_AHBoOo0I,
input
CORETSE_AHBiOo0I,
input
[
7
:
0
]
CORETSE_AHBOIo0I,
input
[
7
:
0
]
CORETSE_AHBIIo0I,
input
CORETSE_AHBlIo0I,
input
[
1
:
0
]
CORETSE_AHBoIo0I,
input
CORETSE_AHBiIo0I,
input
CORETSE_AHBOlo0I,
output
[
15
:
0
]
CORETSE_AHBIlo0I,
output
[
79
:
0
]
CORETSE_AHBllo0I,
output
[
3
:
0
]
CORETSE_AHBolo0I,
output
CORETSE_AHBilo0I
)
;
reg
[
15
:
0
]
CORETSE_AHBO0o0I
;
wire
[
15
:
0
]
CORETSE_AHBI0o0I
;
reg
[
15
:
0
]
CORETSE_AHBl0o0I
;
wire
[
15
:
0
]
CORETSE_AHBo0o0I
;
wire
[
5
:
0
]
CORETSE_AHBi0o0I
;
reg
[
3
:
0
]
CORETSE_AHBO1o0I
;
wire
[
3
:
0
]
CORETSE_AHBI1o0I
;
wire
CORETSE_AHBl1o0I
;
wire
CORETSE_AHBo1o0I
;
reg
CORETSE_AHBi1o0I
;
wire
CORETSE_AHBOoo0I
;
reg
[
7
:
0
]
msg_qu [11 : 0]
;
wire
[
7
:
0
]
msg_qu_c [11 : 0]
;
reg
CORETSE_AHBIoo0I
;
wire
CORETSE_AHBloo0I
;
reg
CORETSE_AHBooo0I
;
reg
CORETSE_AHBioo0I
;
reg
CORETSE_AHBOio0I
;
reg
CORETSE_AHBIio0I
;
reg
CORETSE_AHBlio0I
;
reg
CORETSE_AHBoio0I
;
wire
CORETSE_AHBiio0I
;
reg
CORETSE_AHBOOi0I
;
wire
CORETSE_AHBIOi0I
;
reg
CORETSE_AHBlOi0I
;
wire
CORETSE_AHBoOi0I
;
reg
CORETSE_AHBiOi0I
;
wire
CORETSE_AHBOIi0I
;
reg
CORETSE_AHBIIi0I
;
wire
CORETSE_AHBlIi0I
;
reg
CORETSE_AHBoIi0I
;
wire
CORETSE_AHBiIi0I
;
reg
CORETSE_AHBOli0I
;
wire
CORETSE_AHBIli0I
;
reg
CORETSE_AHBlli0I
;
wire
CORETSE_AHBoli0I
;
reg
CORETSE_AHBili0I
;
wire
CORETSE_AHBO0i0I
;
reg
CORETSE_AHBI0i0I
;
wire
CORETSE_AHBl0i0I
;
reg
CORETSE_AHBo0i0I
;
wire
CORETSE_AHBi0i0I
;
reg
CORETSE_AHBO1i0I
;
wire
CORETSE_AHBI1i0I
;
reg
CORETSE_AHBl1i0I
;
wire
CORETSE_AHBo1i0I
;
reg
CORETSE_AHBi1i0I
;
wire
CORETSE_AHBOoi0I
;
reg
CORETSE_AHBIoi0I
;
wire
CORETSE_AHBloi0I
;
wire
CORETSE_AHBooi0I
;
wire
CORETSE_AHBioi0I
;
wire
CORETSE_AHBOii0I
;
reg
CORETSE_AHBIii0I
;
wire
CORETSE_AHBlii0I
;
reg
CORETSE_AHBoii0I
;
reg
CORETSE_AHBiii0I
;
wire
CORETSE_AHBOOO1I
;
reg
CORETSE_AHBIOO1I
;
wire
CORETSE_AHBlOO1I
;
wire
CORETSE_AHBoOO1I
;
reg
CORETSE_AHBiOO1I
;
wire
CORETSE_AHBOIO1I
;
reg
CORETSE_AHBIIO1I
;
reg
CORETSE_AHBlIO1I
;
wire
CORETSE_AHBoIO1I
;
reg
CORETSE_AHBiIO1I
;
reg
CORETSE_AHBOlO1I
;
reg
[
7
:
0
]
CORETSE_AHBIlO1I
;
wire
[
7
:
0
]
CORETSE_AHBOii0
;
assign
CORETSE_AHBolo0I
=
CORETSE_AHBO1o0I
;
assign
CORETSE_AHBilo0I
=
CORETSE_AHBoio0I
;
assign
CORETSE_AHBllo0I
=
{
msg_qu
[
11
]
,
msg_qu
[
10
]
,
msg_qu
[
9
]
,
msg_qu
[
8
]
,
msg_qu
[
7
]
,
msg_qu
[
6
]
,
msg_qu
[
5
]
,
msg_qu
[
4
]
,
msg_qu
[
3
]
,
msg_qu
[
2
]
}
;
assign
CORETSE_AHBIlo0I
=
{
msg_qu
[
1
]
,
msg_qu
[
0
]
}
;
assign
CORETSE_AHBOii0
=
{
8
{
CORETSE_AHBoIo0I
[
1
]
}
}
&
CORETSE_AHBOIo0I
|
{
8
{
~
CORETSE_AHBoIo0I
[
1
]
}
}
&
CORETSE_AHBIlO1I
;
assign
CORETSE_AHBOOO1I
=
~
CORETSE_AHBIii0I
&
CORETSE_AHBlIo0I
;
assign
CORETSE_AHBoOO1I
=
CORETSE_AHBOOO1I
|
CORETSE_AHBIOO1I
;
assign
CORETSE_AHBlOO1I
=
CORETSE_AHBoIo0I
[
1
]
&
CORETSE_AHBOOO1I
|
~
CORETSE_AHBoIo0I
[
1
]
&
CORETSE_AHBiOO1I
;
assign
CORETSE_AHBOIO1I
=
CORETSE_AHBoIo0I
[
1
]
|
~
CORETSE_AHBoIo0I
[
1
]
&
(
CORETSE_AHBlIO1I
&
~
CORETSE_AHBIIO1I
)
;
assign
CORETSE_AHBoIO1I
=
~
CORETSE_AHBOlO1I
&
(
CORETSE_AHBOOO1I
|
(
~
CORETSE_AHBOOO1I
&
CORETSE_AHBlIO1I
)
)
;
assign
CORETSE_AHBlii0I
=
CORETSE_AHBIOo0I
|
CORETSE_AHBlOo0I
;
assign
CORETSE_AHBi0o0I
=
{
CORETSE_AHBOii0
[
3
:
0
]
,
2
'b
00
}
-
2
'b
10
;
assign
CORETSE_AHBiio0I
=
~
CORETSE_AHBIio0I
&
(
CORETSE_AHBIoo0I
|
(
~
CORETSE_AHBIoo0I
&
CORETSE_AHBlio0I
)
)
;
assign
CORETSE_AHBIOi0I
=
CORETSE_AHBiIo0I
|
(
CORETSE_AHBOOi0I
&
~
(
CORETSE_AHBioo0I
&
CORETSE_AHBlOO1I
)
|
CORETSE_AHBlli0I
&
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
8
&&
CORETSE_AHBOii0
!=
8
'h
11
)
|
CORETSE_AHBili0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
&&
CORETSE_AHBOii0
!=
8
'h
11
)
|
CORETSE_AHBi1i0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
2
&&
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
!=
16
'h
013F
)
|
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
0
)
&
(
CORETSE_AHBIIo0I
[
3
]
==
1
'b
1
)
|
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
1F
)
|
(
!
CORETSE_AHBoOi0I
&
!
CORETSE_AHBOIi0I
&
!
CORETSE_AHBlIi0I
&
!
CORETSE_AHBiIi0I
&
!
CORETSE_AHBIli0I
&
!
CORETSE_AHBoli0I
&
!
CORETSE_AHBO0i0I
&
!
CORETSE_AHBl0i0I
&
!
CORETSE_AHBi0i0I
&
!
CORETSE_AHBI1i0I
&
!
CORETSE_AHBo1i0I
&
!
CORETSE_AHBOoi0I
&
!
CORETSE_AHBloi0I
)
)
;
assign
CORETSE_AHBoOi0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBOOi0I
&
CORETSE_AHBioo0I
&
CORETSE_AHBlOO1I
&
CORETSE_AHBlIo0I
|
CORETSE_AHBlOi0I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
A
)
)
;
assign
CORETSE_AHBOIi0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBlOi0I
&
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
A
)
)
;
assign
CORETSE_AHBlIi0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBiOi0I
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
8100
)
|
CORETSE_AHBoIi0I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
8100
)
|
CORETSE_AHBIIi0I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
;
assign
CORETSE_AHBiIi0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBiOi0I
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
88A8
)
|
CORETSE_AHBoIi0I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
88A8
)
|
CORETSE_AHBoIi0I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
;
assign
CORETSE_AHBIli0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBiOi0I
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
8847
||
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
8848
)
|
CORETSE_AHBIIi0I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
8847
||
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
8848
)
|
CORETSE_AHBOli0I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
;
assign
CORETSE_AHBoli0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBOli0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
&
(
CORETSE_AHBOii0
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBOii0
[
3
:
0
]
>
4
'h
4
)
|
CORETSE_AHBI0i0I
&
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
&
(
CORETSE_AHBOii0
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBOii0
[
3
:
0
]
>
4
'h
4
)
|
CORETSE_AHBlli0I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
8
&&
CORETSE_AHBOii0
!=
8
'h
11
)
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
;
assign
CORETSE_AHBO0i0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBOli0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
&
(
CORETSE_AHBOii0
[
7
:
4
]
==
4
'h
6
)
|
CORETSE_AHBo0i0I
&
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
|
CORETSE_AHBili0I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
;
assign
CORETSE_AHBl0i0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBiOi0I
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
0800
)
|
CORETSE_AHBIIi0I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
0800
)
|
CORETSE_AHBI0i0I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
;
assign
CORETSE_AHBi0i0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBiOi0I
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
86DD
)
|
CORETSE_AHBIIi0I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
86DD
)
|
CORETSE_AHBo0i0I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
;
assign
CORETSE_AHBI1i0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBiOi0I
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
88F7
)
|
CORETSE_AHBIIi0I
&
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
&
(
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
==
16
'h
88F7
)
)
;
assign
CORETSE_AHBo1i0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBili0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
&&
CORETSE_AHBOii0
==
8
'h
11
)
|
CORETSE_AHBl1i0I
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
;
assign
CORETSE_AHBOoi0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBlli0I
&
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
|
CORETSE_AHBl1i0I
&
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
|
CORETSE_AHBi1i0I
&
~
(
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
2
&&
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
!=
16
'h
013F
)
)
&
~
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
)
;
assign
CORETSE_AHBloi0I
=
~
CORETSE_AHBiIo0I
&
(
CORETSE_AHBO1i0I
|
CORETSE_AHBi1i0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
|
CORETSE_AHBIoi0I
&
!
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
1F
)
&
!
(
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
0
)
&
(
(
CORETSE_AHBOii0
[
2
]
|
CORETSE_AHBOii0
[
3
]
)
==
1
'b
1
)
)
)
;
assign
CORETSE_AHBI1o0I
=
{
4
{
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
0
)
}
}
&
CORETSE_AHBOii0
[
3
:
0
]
|
{
4
{
~
(
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
0
)
)
}
}
&
CORETSE_AHBO1o0I
;
assign
CORETSE_AHBloo0I
=
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
1F
)
;
assign
CORETSE_AHBl1o0I
=
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
13
)
;
assign
CORETSE_AHBo1o0I
=
CORETSE_AHBIoi0I
&
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
1F
)
;
assign
CORETSE_AHBI0o0I
=
{
16
{
(
CORETSE_AHBlOi0I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
A
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBoIi0I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBIIi0I
&
!
(
CORETSE_AHBO0o0I
[
1
:
0
]
==
2
'h
3
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBOli0I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBI0i0I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBo0i0I
&
!
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBl1i0I
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBlli0I
&
!
(
CORETSE_AHBO0o0I
[
3
:
0
]
==
4
'h
8
&&
CORETSE_AHBOii0
!=
8
'h
11
)
&
!
(
CORETSE_AHBO0o0I
==
CORETSE_AHBl0o0I
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBili0I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBi1i0I
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
2
&&
{
CORETSE_AHBOii0
,
CORETSE_AHBIIo0I
}
!=
16
'h
013F
)
&
!
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
7
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
|
{
16
{
(
CORETSE_AHBIoi0I
&
!
(
CORETSE_AHBO0o0I
[
4
:
0
]
==
5
'h
1F
)
)
}
}
&
(
CORETSE_AHBO0o0I
+
1
'b
1
)
;
assign
CORETSE_AHBooi0I
=
CORETSE_AHBOli0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
5
)
&
(
CORETSE_AHBOii0
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBOii0
[
3
:
0
]
>
4
'h
4
)
;
assign
CORETSE_AHBioi0I
=
CORETSE_AHBI0i0I
&
(
CORETSE_AHBO0o0I
[
0
]
==
1
'h
1
)
&
(
CORETSE_AHBOii0
[
7
:
4
]
==
4
'h
4
&&
CORETSE_AHBOii0
[
3
:
0
]
>
4
'h
4
)
;
assign
CORETSE_AHBOii0I
=
CORETSE_AHBili0I
&
(
CORETSE_AHBO0o0I
[
2
:
0
]
==
3
'h
3
)
;
assign
CORETSE_AHBo0o0I
=
{
16
{
CORETSE_AHBooi0I
}
}
&
{
10
'b
0
,
CORETSE_AHBi0o0I
}
|
{
16
{
CORETSE_AHBioi0I
}
}
&
{
10
'b
0
,
CORETSE_AHBi0o0I
}
|
{
16
{
CORETSE_AHBOii0I
}
}
&
(
16
'h
28
-
16
'h
8
)
|
{
16
{
~
(
CORETSE_AHBooi0I
|
CORETSE_AHBioi0I
|
CORETSE_AHBOii0I
)
}
}
&
CORETSE_AHBl0o0I
;
assign
CORETSE_AHBOoo0I
=
~
CORETSE_AHBo1o0I
&
(
CORETSE_AHBl1o0I
|
(
~
CORETSE_AHBl1o0I
&
CORETSE_AHBi1o0I
)
)
;
assign
msg_qu_c
[
0
]
=
(
{
8
{
CORETSE_AHBi1o0I
}
}
&
CORETSE_AHBOii0
)
|
(
{
8
{
~
CORETSE_AHBi1o0I
}
}
&
msg_qu
[
0
]
)
;
generate
genvar
CORETSE_AHBOloI
;
for
(
CORETSE_AHBOloI
=
1
;
CORETSE_AHBOloI
<
12
;
CORETSE_AHBOloI
=
CORETSE_AHBOloI
+
1
)
begin
:
CORETSE_AHBllO1I
assign
msg_qu_c
[
CORETSE_AHBOloI
]
=
(
{
8
{
CORETSE_AHBi1o0I
}
}
&
msg_qu
[
CORETSE_AHBOloI
-
1
]
)
|
(
{
8
{
~
CORETSE_AHBi1o0I
}
}
&
msg_qu
[
CORETSE_AHBOloI
]
)
;
end
endgenerate
always
@
(
posedge
CORETSE_AHBOOo0I
or
posedge
CORETSE_AHBiii0I
)
begin
if
(
CORETSE_AHBiii0I
)
begin
CORETSE_AHBooo0I
<=
1
'b
0
;
CORETSE_AHBioo0I
<=
1
'b
0
;
CORETSE_AHBOio0I
<=
1
'b
0
;
CORETSE_AHBIio0I
<=
1
'b
0
;
CORETSE_AHBO0o0I
<=
16
'b
0
;
CORETSE_AHBl0o0I
<=
16
'b
0
;
CORETSE_AHBO1o0I
<=
4
'b
0
;
CORETSE_AHBi1o0I
<=
1
'b
0
;
msg_qu
[
0
]
<=
8
'b
0
;
msg_qu
[
1
]
<=
8
'b
0
;
msg_qu
[
2
]
<=
8
'b
0
;
msg_qu
[
3
]
<=
8
'b
0
;
msg_qu
[
4
]
<=
8
'b
0
;
msg_qu
[
5
]
<=
8
'b
0
;
msg_qu
[
6
]
<=
8
'b
0
;
msg_qu
[
7
]
<=
8
'b
0
;
msg_qu
[
8
]
<=
8
'b
0
;
msg_qu
[
9
]
<=
8
'b
0
;
msg_qu
[
10
]
<=
8
'b
0
;
msg_qu
[
11
]
<=
8
'b
0
;
CORETSE_AHBIoo0I
<=
1
'b
0
;
CORETSE_AHBlio0I
<=
1
'b
0
;
CORETSE_AHBoio0I
<=
1
'b
0
;
CORETSE_AHBOOi0I
<=
1
'b
1
;
CORETSE_AHBlOi0I
<=
1
'b
0
;
CORETSE_AHBiOi0I
<=
1
'b
0
;
CORETSE_AHBIIi0I
<=
1
'b
0
;
CORETSE_AHBoIi0I
<=
1
'b
0
;
CORETSE_AHBOli0I
<=
1
'b
0
;
CORETSE_AHBlli0I
<=
1
'b
0
;
CORETSE_AHBili0I
<=
1
'b
0
;
CORETSE_AHBI0i0I
<=
1
'b
0
;
CORETSE_AHBo0i0I
<=
1
'b
0
;
CORETSE_AHBO1i0I
<=
1
'b
0
;
CORETSE_AHBl1i0I
<=
1
'b
0
;
CORETSE_AHBi1i0I
<=
1
'b
0
;
CORETSE_AHBIoi0I
<=
1
'b
0
;
CORETSE_AHBIii0I
<=
1
'b
0
;
CORETSE_AHBIOO1I
<=
1
'b
0
;
CORETSE_AHBiOO1I
<=
1
'b
0
;
CORETSE_AHBIIO1I
<=
1
'b
0
;
CORETSE_AHBlIO1I
<=
1
'b
0
;
CORETSE_AHBiIO1I
<=
1
'b
0
;
CORETSE_AHBOlO1I
<=
1
'b
0
;
CORETSE_AHBIlO1I
<=
8
'b
0
;
end
else
begin
CORETSE_AHBooo0I
<=
CORETSE_AHBoOo0I
;
CORETSE_AHBioo0I
<=
CORETSE_AHBooo0I
;
CORETSE_AHBOio0I
<=
CORETSE_AHBOlo0I
;
CORETSE_AHBIio0I
<=
CORETSE_AHBOio0I
;
CORETSE_AHBlio0I
<=
CORETSE_AHBiio0I
;
CORETSE_AHBoio0I
<=
CORETSE_AHBlio0I
;
CORETSE_AHBIii0I
<=
CORETSE_AHBlIo0I
;
CORETSE_AHBIOO1I
<=
CORETSE_AHBOOO1I
;
CORETSE_AHBiOO1I
<=
CORETSE_AHBoOO1I
;
CORETSE_AHBIIO1I
<=
CORETSE_AHBOIO1I
;
CORETSE_AHBlIO1I
<=
CORETSE_AHBoIO1I
;
CORETSE_AHBiIO1I
<=
CORETSE_AHBiIo0I
;
CORETSE_AHBOlO1I
<=
CORETSE_AHBiIO1I
;
CORETSE_AHBIlO1I
<=
CORETSE_AHBOIo0I
;
if
(
CORETSE_AHBiOo0I
&&
CORETSE_AHBIIO1I
)
begin
CORETSE_AHBO0o0I
<=
CORETSE_AHBI0o0I
;
CORETSE_AHBl0o0I
<=
CORETSE_AHBo0o0I
;
CORETSE_AHBO1o0I
<=
CORETSE_AHBI1o0I
;
CORETSE_AHBi1o0I
<=
CORETSE_AHBOoo0I
;
msg_qu
[
0
]
<=
msg_qu_c
[
0
]
;
msg_qu
[
1
]
<=
msg_qu_c
[
1
]
;
msg_qu
[
2
]
<=
msg_qu_c
[
2
]
;
msg_qu
[
3
]
<=
msg_qu_c
[
3
]
;
msg_qu
[
4
]
<=
msg_qu_c
[
4
]
;
msg_qu
[
5
]
<=
msg_qu_c
[
5
]
;
msg_qu
[
6
]
<=
msg_qu_c
[
6
]
;
msg_qu
[
7
]
<=
msg_qu_c
[
7
]
;
msg_qu
[
8
]
<=
msg_qu_c
[
8
]
;
msg_qu
[
9
]
<=
msg_qu_c
[
9
]
;
msg_qu
[
10
]
<=
msg_qu_c
[
10
]
;
msg_qu
[
11
]
<=
msg_qu_c
[
11
]
;
CORETSE_AHBIoo0I
<=
CORETSE_AHBloo0I
;
CORETSE_AHBOOi0I
<=
CORETSE_AHBIOi0I
;
CORETSE_AHBlOi0I
<=
CORETSE_AHBoOi0I
;
CORETSE_AHBiOi0I
<=
CORETSE_AHBOIi0I
;
CORETSE_AHBIIi0I
<=
CORETSE_AHBlIi0I
;
CORETSE_AHBoIi0I
<=
CORETSE_AHBiIi0I
;
CORETSE_AHBOli0I
<=
CORETSE_AHBIli0I
;
CORETSE_AHBlli0I
<=
CORETSE_AHBoli0I
;
CORETSE_AHBili0I
<=
CORETSE_AHBO0i0I
;
CORETSE_AHBI0i0I
<=
CORETSE_AHBl0i0I
;
CORETSE_AHBo0i0I
<=
CORETSE_AHBi0i0I
;
CORETSE_AHBO1i0I
<=
CORETSE_AHBI1i0I
;
CORETSE_AHBl1i0I
<=
CORETSE_AHBo1i0I
;
CORETSE_AHBi1i0I
<=
CORETSE_AHBOoi0I
;
CORETSE_AHBIoi0I
<=
CORETSE_AHBloi0I
;
end
end
end
always
@
(
posedge
CORETSE_AHBOOo0I
or
posedge
CORETSE_AHBlii0I
)
begin
if
(
CORETSE_AHBlii0I
)
begin
CORETSE_AHBoii0I
<=
1
'b
1
;
CORETSE_AHBiii0I
<=
1
'b
1
;
end
else
begin
CORETSE_AHBoii0I
<=
1
'b
0
;
CORETSE_AHBiii0I
<=
CORETSE_AHBoii0I
;
end
end
endmodule
