// REVISION    : $Revision: 1.12 $
//         Mentor Graphics Corporation Proprietary and Confidential
//         Copyright Mentor Graphics Corporation and Licensors 2004
`include "include.v"
module
slave
(
HWDATA
,
HADDR
,
HSEL
,
HTRANS
,
HWRITE
,
HCLK
,
CORETSE_AHBl1Il
,
HRDATA
,
HRESP
,
HREADY
,
CORETSE_AHBIil0
,
CORETSE_AHBioOl
,
CORETSE_AHBIoll
,
CORETSE_AHBlIIl
,
CORETSE_AHBOiOl
,
CORETSE_AHBloll
,
CORETSE_AHBIiOl
,
CORETSE_AHBliOl
,
CORETSE_AHBi0l0
,
CORETSE_AHBO1l0
)
;
input
[
31
:
0
]
HWDATA
;
input
[
9
:
2
]
HADDR
;
input
HSEL
;
input
[
1
:
0
]
HTRANS
;
input
HWRITE
;
input
HREADY
;
input
HCLK
;
input
CORETSE_AHBl1Il
;
output
[
31
:
0
]
HRDATA
;
output
[
1
:
0
]
HRESP
;
output
CORETSE_AHBIil0
;
output
CORETSE_AHBioOl
;
output
CORETSE_AHBIoll
;
output
CORETSE_AHBlIIl
;
output
[
7
:
0
]
CORETSE_AHBOiOl
;
output
[
31
:
0
]
CORETSE_AHBloll
;
input
[
31
:
0
]
CORETSE_AHBIiOl
;
input
CORETSE_AHBliOl
;
output
CORETSE_AHBi0l0
;
input
CORETSE_AHBO1l0
;
reg
CORETSE_AHBioOl
;
reg
CORETSE_AHBIoll
;
reg
CORETSE_AHBlIIl
;
reg
[
7
:
0
]
CORETSE_AHBOiOl
;
reg
CORETSE_AHBoI0oI
;
reg
[
31
:
0
]
CORETSE_AHBiI0oI
;
reg
[
2
:
0
]
CORETSE_AHBOl0oI
;
reg
CORETSE_AHBIl0oI
;
reg
CORETSE_AHBll0oI
;
reg
CORETSE_AHBi0l0
;
wire
[
1
:
0
]
HRESP
;
wire
CORETSE_AHBol0oI
;
wire
CORETSE_AHBil0oI
;
assign
CORETSE_AHBil0oI
=
~
HADDR
[
9
]
&
(
HADDR
[
8
]
^
HADDR
[
7
]
)
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBO00oI
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBoI0oI
<=
1
;
CORETSE_AHBioOl
<=
1
;
CORETSE_AHBOiOl
<=
0
;
CORETSE_AHBIoll
<=
1
;
CORETSE_AHBlIIl
<=
1
;
end
else
begin
if
(
HREADY
)
begin
CORETSE_AHBioOl
<=
!
(
HSEL
&&
(
(
HTRANS
==
`CORETSE_AHBIi1l
)
||
(
HTRANS
==
`CORETSE_AHBoi1l
)
)
&&
!
CORETSE_AHBil0oI
)
;
CORETSE_AHBlIIl
<=
!
(
HSEL
&&
(
(
HTRANS
==
`CORETSE_AHBIi1l
)
||
(
HTRANS
==
`CORETSE_AHBoi1l
)
)
&&
CORETSE_AHBil0oI
)
;
CORETSE_AHBOiOl
<=
HADDR
;
CORETSE_AHBIoll
<=
!
HWRITE
;
end
CORETSE_AHBoI0oI
<=
CORETSE_AHBol0oI
;
end
end
assign
CORETSE_AHBol0oI
=
!
CORETSE_AHBIoll
||
CORETSE_AHBioOl
||
CORETSE_AHBliOl
;
assign
CORETSE_AHBIil0
=
CORETSE_AHBIl0oI
?
CORETSE_AHBll0oI
:
!
(
!
CORETSE_AHBol0oI
&&
CORETSE_AHBoI0oI
)
;
assign
HRESP
=
(
!
CORETSE_AHBol0oI
)
?
`CORETSE_AHBI1il
:
`CORETSE_AHBiool
;
assign
CORETSE_AHBloll
=
HWDATA
;
assign
HRDATA
=
CORETSE_AHBIl0oI
?
CORETSE_AHBiI0oI
:
CORETSE_AHBIiOl
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBI00oI
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBIl0oI
<=
0
;
CORETSE_AHBll0oI
<=
0
;
CORETSE_AHBi0l0
<=
0
;
CORETSE_AHBOl0oI
<=
0
;
CORETSE_AHBiI0oI
<=
0
;
end
else
begin
CORETSE_AHBOl0oI
<=
{
CORETSE_AHBOl0oI
[
1
:
0
]
,
CORETSE_AHBO1l0
}
;
if
(
HREADY
)
begin
CORETSE_AHBIl0oI
<=
HSEL
&&
CORETSE_AHBil0oI
&&
(
(
HTRANS
==
`CORETSE_AHBIi1l
)
||
(
HTRANS
==
`CORETSE_AHBoi1l
)
)
;
CORETSE_AHBll0oI
<=
0
;
CORETSE_AHBi0l0
<=
HSEL
&&
CORETSE_AHBil0oI
&&
(
(
HTRANS
==
`CORETSE_AHBIi1l
)
||
(
HTRANS
==
`CORETSE_AHBoi1l
)
)
&&
!
CORETSE_AHBOl0oI
[
1
]
;
end
else
if
(
CORETSE_AHBIl0oI
)
CORETSE_AHBi0l0
<=
!
CORETSE_AHBOl0oI
[
1
]
;
if
(
CORETSE_AHBOl0oI
[
2
:
1
]
==
2
'b
01
)
begin
CORETSE_AHBi0l0
<=
0
;
CORETSE_AHBiI0oI
<=
CORETSE_AHBIiOl
;
CORETSE_AHBll0oI
<=
1
;
end
end
end
endmodule
