// REVISION    : $Revision: 1.1 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
pecar
(
CORETSE_AHBO111
,
CORETSE_AHBI111
,
CORETSE_AHBl111
,
CORETSE_AHBiOO1
,
CORETSE_AHBo1Oo
,
CORETSE_AHBoi0
,
CORETSE_AHBllo
,
CORETSE_AHBo111
,
CORETSE_AHBi1Oo
,
CORETSE_AHBii0
,
CORETSE_AHBl0o
,
CORETSE_AHBio11
,
CORETSE_AHBoOIo
,
CORETSE_AHBiOIo
,
CORETSE_AHBo011
,
CORETSE_AHBOi1
,
CORETSE_AHBio1
,
CORETSE_AHBii01
,
CORETSE_AHBllOo
,
CORETSE_AHBolOo
,
CORETSE_AHBilOo
,
CORETSE_AHBO0Oo
,
CORETSE_AHBI0Oo
,
CORETSE_AHBOIIo
,
CORETSE_AHBIIIo
,
CORETSE_AHBl0Oo
,
CORETSE_AHBOOIo
,
CORETSE_AHBIOIo
,
CORETSE_AHBoo1
,
CORETSE_AHBIi11
,
CORETSE_AHBli11
,
CORETSE_AHBoi11
,
CORETSE_AHBii11
,
CORETSE_AHBoio1
,
CORETSE_AHBiio1
,
CORETSE_AHBIio1
,
CORETSE_AHBlio1
,
CORETSE_AHBo0Oo
,
CORETSE_AHBi0Oo
,
CORETSE_AHBII11
,
CORETSE_AHBoI11
,
CORETSE_AHBO1Oo
,
CORETSE_AHBllo1
,
CORETSE_AHBolo1
,
CORETSE_AHBilo1
,
CORETSE_AHBlIIo
,
CORETSE_AHBoIIo
,
CORETSE_AHBiIIo
)
;
input
CORETSE_AHBO111
,
CORETSE_AHBI111
,
CORETSE_AHBl111
;
input
CORETSE_AHBiOO1
,
CORETSE_AHBo1Oo
;
input
CORETSE_AHBoi0
,
CORETSE_AHBllo
;
input
CORETSE_AHBo111
,
CORETSE_AHBi1Oo
;
input
CORETSE_AHBii0
,
CORETSE_AHBl0o
;
input
CORETSE_AHBio11
;
input
CORETSE_AHBoOIo
,
CORETSE_AHBiOIo
,
CORETSE_AHBo011
;
input
CORETSE_AHBOi1
,
CORETSE_AHBio1
,
CORETSE_AHBii01
;
input
CORETSE_AHBllOo
,
CORETSE_AHBolOo
,
CORETSE_AHBilOo
,
CORETSE_AHBO0Oo
;
input
CORETSE_AHBI0Oo
,
CORETSE_AHBOIIo
,
CORETSE_AHBIIIo
;
input
CORETSE_AHBl0Oo
;
input
CORETSE_AHBOOIo
,
CORETSE_AHBIOIo
;
input
CORETSE_AHBoo1
;
output
CORETSE_AHBIi11
,
CORETSE_AHBli11
;
output
CORETSE_AHBoi11
,
CORETSE_AHBii11
;
output
CORETSE_AHBoio1
,
CORETSE_AHBiio1
;
output
CORETSE_AHBIio1
,
CORETSE_AHBlio1
,
CORETSE_AHBo0Oo
,
CORETSE_AHBi0Oo
;
output
CORETSE_AHBII11
,
CORETSE_AHBoI11
;
output
CORETSE_AHBO1Oo
;
output
CORETSE_AHBllo1
;
output
CORETSE_AHBolo1
;
output
CORETSE_AHBilo1
;
output
CORETSE_AHBlIIo
;
output
CORETSE_AHBoIIo
;
output
CORETSE_AHBiIIo
;
parameter
CORETSE_AHBIoII
=
1
;
wire
CORETSE_AHBi0lo
;
reg
CORETSE_AHBO1lo
,
CORETSE_AHBI1lo
;
wire
CORETSE_AHBl1lo
;
wire
CORETSE_AHBo1lo
;
reg
CORETSE_AHBi1lo
,
CORETSE_AHBOolo
;
wire
CORETSE_AHBIolo
;
wire
CORETSE_AHBlolo
;
reg
CORETSE_AHBoolo
,
CORETSE_AHBiolo
;
wire
CORETSE_AHBOilo
;
wire
CORETSE_AHBIilo
;
reg
CORETSE_AHBlilo
,
CORETSE_AHBoilo
;
wire
CORETSE_AHBiilo
;
wire
CORETSE_AHBOO0o
;
reg
CORETSE_AHBIO0o
,
CORETSE_AHBlO0o
;
wire
CORETSE_AHBoO0o
;
wire
CORETSE_AHBiO0o
;
reg
CORETSE_AHBOI0o
,
CORETSE_AHBII0o
;
wire
CORETSE_AHBlI0o
;
wire
CORETSE_AHBoI0o
;
reg
CORETSE_AHBiI0o
,
CORETSE_AHBOl0o
;
wire
CORETSE_AHBIl0o
;
wire
CORETSE_AHBll0o
;
reg
CORETSE_AHBol0o
,
CORETSE_AHBil0o
;
wire
CORETSE_AHBO00o
;
wire
CORETSE_AHBI00o
;
reg
CORETSE_AHBl00o
,
CORETSE_AHBo00o
;
wire
CORETSE_AHBi00o
;
reg
CORETSE_AHBO10o
,
CORETSE_AHBI10o
;
wire
CORETSE_AHBl10o
;
reg
CORETSE_AHBo10o
;
reg
CORETSE_AHBi10o
;
wire
CORETSE_AHBOo0o
;
wire
CORETSE_AHBIo0o
;
reg
CORETSE_AHBlo0o
,
CORETSE_AHBoo0o
;
wire
CORETSE_AHBio0o
;
reg
CORETSE_AHBOi0o
,
CORETSE_AHBIi0o
;
wire
CORETSE_AHBli0o
;
reg
CORETSE_AHBoi0o
,
CORETSE_AHBii0o
;
wire
CORETSE_AHBOO1o
;
wire
CORETSE_AHBIO1o
;
reg
CORETSE_AHBlO1o
,
CORETSE_AHBoO1o
;
wire
CORETSE_AHBiO1o
;
reg
CORETSE_AHBOI1o
,
CORETSE_AHBII1o
;
wire
CORETSE_AHBlI1o
;
wire
CORETSE_AHBoI1o
;
wire
CORETSE_AHBiI1o
;
assign
CORETSE_AHBi0lo
=
CORETSE_AHBio1
|
CORETSE_AHBii01
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBO1lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0lo
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBI1lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1lo
;
end
assign
CORETSE_AHBl1lo
=
CORETSE_AHBi0lo
|
CORETSE_AHBI1lo
;
assign
CORETSE_AHBoio1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBl1lo
;
assign
CORETSE_AHBo1lo
=
CORETSE_AHBio1
|
CORETSE_AHBii01
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBi1lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1lo
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBOolo
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1lo
;
end
assign
CORETSE_AHBIolo
=
CORETSE_AHBo1lo
|
CORETSE_AHBOolo
;
assign
CORETSE_AHBiio1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBIolo
;
assign
CORETSE_AHBlolo
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBllOo
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBoolo
<=
#
CORETSE_AHBIoII
CORETSE_AHBlolo
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBiolo
<=
#
CORETSE_AHBIoII
CORETSE_AHBoolo
;
end
assign
CORETSE_AHBOilo
=
CORETSE_AHBlolo
|
CORETSE_AHBiolo
;
assign
CORETSE_AHBIio1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBOilo
;
assign
CORETSE_AHBIilo
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBolOo
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBlilo
<=
#
CORETSE_AHBIoII
CORETSE_AHBIilo
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBoilo
<=
#
CORETSE_AHBIoII
CORETSE_AHBlilo
;
end
assign
CORETSE_AHBiilo
=
CORETSE_AHBIilo
|
CORETSE_AHBoilo
;
assign
CORETSE_AHBlio1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBiilo
;
assign
CORETSE_AHBOO0o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBOIIo
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBIO0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBOO0o
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBlO0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIO0o
;
end
assign
CORETSE_AHBoO0o
=
CORETSE_AHBOO0o
|
CORETSE_AHBlO0o
;
assign
CORETSE_AHBII11
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBoO0o
;
assign
CORETSE_AHBiO0o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBIIIo
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBOI0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO0o
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBII0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBOI0o
;
end
assign
CORETSE_AHBlI0o
=
CORETSE_AHBiO0o
|
CORETSE_AHBII0o
;
assign
CORETSE_AHBoI11
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBlI0o
;
assign
CORETSE_AHBoI0o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBilOo
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBiI0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI0o
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBOl0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBiI0o
;
end
assign
CORETSE_AHBIl0o
=
CORETSE_AHBoI0o
|
CORETSE_AHBOl0o
;
assign
CORETSE_AHBo0Oo
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBIl0o
;
assign
CORETSE_AHBll0o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBO0Oo
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBol0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBll0o
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBil0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0o
;
end
assign
CORETSE_AHBO00o
=
CORETSE_AHBll0o
|
CORETSE_AHBil0o
;
assign
CORETSE_AHBi0Oo
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBO00o
;
assign
CORETSE_AHBI00o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBI0Oo
;
always
@
(
posedge
CORETSE_AHBio11
)
begin
CORETSE_AHBl00o
<=
#
CORETSE_AHBIoII
CORETSE_AHBI00o
;
end
always
@
(
posedge
CORETSE_AHBio11
)
begin
CORETSE_AHBo00o
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00o
;
end
assign
CORETSE_AHBi00o
=
CORETSE_AHBI00o
|
CORETSE_AHBo00o
;
assign
CORETSE_AHBO1Oo
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBi00o
;
always
@
(
posedge
CORETSE_AHBO111
)
begin
CORETSE_AHBO10o
<=
#
CORETSE_AHBIoII
CORETSE_AHBio1
;
end
always
@
(
posedge
CORETSE_AHBO111
)
begin
CORETSE_AHBI10o
<=
#
CORETSE_AHBIoII
CORETSE_AHBO10o
;
end
assign
CORETSE_AHBl10o
=
CORETSE_AHBio1
|
CORETSE_AHBI10o
;
always
@
(
posedge
CORETSE_AHBO111
)
begin
if
(
CORETSE_AHBl10o
)
CORETSE_AHBo10o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo10o
<=
#
CORETSE_AHBIoII
~
CORETSE_AHBo10o
;
end
assign
CORETSE_AHBIi11
=
(
CORETSE_AHBl111
)
?
CORETSE_AHBo10o
:
CORETSE_AHBiOO1
;
assign
CORETSE_AHBli11
=
CORETSE_AHBo1Oo
;
always
@
(
posedge
CORETSE_AHBO111
)
begin
if
(
CORETSE_AHBl10o
)
CORETSE_AHBi10o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi10o
<=
#
CORETSE_AHBIoII
~
CORETSE_AHBi10o
;
end
assign
CORETSE_AHBOo0o
=
(
CORETSE_AHBl111
)
?
CORETSE_AHBi10o
:
CORETSE_AHBo111
;
assign
CORETSE_AHBoi11
=
(
CORETSE_AHBoo1
|
~
CORETSE_AHBo011
)
&
CORETSE_AHBOo0o
|
(
~
CORETSE_AHBoo1
&
CORETSE_AHBo011
)
&
CORETSE_AHBoOIo
;
assign
CORETSE_AHBii11
=
(
CORETSE_AHBoo1
|
~
CORETSE_AHBo011
)
&
CORETSE_AHBi1Oo
|
(
~
CORETSE_AHBoo1
&
CORETSE_AHBo011
)
&
CORETSE_AHBiOIo
;
assign
CORETSE_AHBIo0o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBl0Oo
;
always
@
(
posedge
CORETSE_AHBI111
)
begin
CORETSE_AHBlo0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo0o
;
end
always
@
(
posedge
CORETSE_AHBI111
)
begin
CORETSE_AHBoo0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo0o
;
end
assign
CORETSE_AHBio0o
=
CORETSE_AHBIo0o
|
CORETSE_AHBoo0o
;
assign
CORETSE_AHBllo1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBio0o
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBOi0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo0o
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBIi0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi0o
;
end
assign
CORETSE_AHBli0o
=
CORETSE_AHBIo0o
|
CORETSE_AHBIi0o
;
assign
CORETSE_AHBolo1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBli0o
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBoi0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo0o
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBii0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBoi0o
;
end
assign
CORETSE_AHBOO1o
=
CORETSE_AHBIo0o
|
CORETSE_AHBii0o
;
assign
CORETSE_AHBilo1
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBOO1o
;
assign
CORETSE_AHBIO1o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBOOIo
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBlO1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIO1o
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBoO1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO1o
;
end
assign
CORETSE_AHBiO1o
=
CORETSE_AHBIO1o
|
CORETSE_AHBoO1o
;
assign
CORETSE_AHBlIIo
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBiO1o
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBOI1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBIO1o
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBII1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBOI1o
;
end
assign
CORETSE_AHBlI1o
=
CORETSE_AHBIO1o
|
CORETSE_AHBII1o
;
assign
CORETSE_AHBoIIo
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBlI1o
;
assign
CORETSE_AHBoI1o
=
CORETSE_AHBio1
|
CORETSE_AHBii01
|
CORETSE_AHBIOIo
;
assign
CORETSE_AHBiI1o
=
CORETSE_AHBoI1o
;
assign
CORETSE_AHBiIIo
=
CORETSE_AHBoo1
?
CORETSE_AHBio1
:
CORETSE_AHBiI1o
;
endmodule
