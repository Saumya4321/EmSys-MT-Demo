//                        Proprietary and Confidential 
// REVISION    : $Revision: 1.57 $ 
module
tsmac_top
#
(
parameter
TABITS
=
12
,
parameter
RABITS
=
12
,
parameter
MCXMAC_SAL_ON
=
0
,
parameter
MCXMAC_WOL_ON
=
0
,
parameter
MCXMAC_STATS_ON
=
0
,
parameter
CORETSE_AHBoOI
=
0
,
parameter
CORETSE_AHBiOI
=
0
,
parameter
CORETSE_AHBlOI
=
0
,
parameter
CORETSE_AHBIII
=
1
,
parameter
CORETSE_AHBlII
=
2
,
parameter
CORETSE_AHBoII
=
1
,
parameter
CORETSE_AHBiII
=
2
,
parameter
CORETSE_AHBOlI
=
18
,
parameter
CORETSE_AHBIlI
=
18
,
parameter
CORETSE_AHBllI
=
5
,
parameter
CORETSE_AHBolI
=
5
,
parameter
CORETSE_AHBOII
=
1
)
(
input
CORETSE_AHBO0I,
input
CORETSE_AHBI0I,
input
CORETSE_AHBl0I,
input
CORETSE_AHBo0I,
input
CORETSE_AHBi0I,
input
CORETSE_AHBO1I,
input
[
7
:
0
]
CORETSE_AHBI1I,
input
CORETSE_AHBl1I,
output
CORETSE_AHBo1I,
output
[
7
:
0
]
CORETSE_AHBi1I,
output
CORETSE_AHBOoI,
input
CORETSE_AHBIoI,
input
CORETSE_AHBloI,
input
[
31
:
0
]
CORETSE_AHBioI,
input
[
9
:
2
]
CORETSE_AHBOiI,
input
CORETSE_AHBIiI,
input
[
1
:
0
]
CORETSE_AHBliI,
input
CORETSE_AHBoiI,
output
[
31
:
0
]
CORETSE_AHBiiI,
output
[
1
:
0
]
CORETSE_AHBOOl,
output
CORETSE_AHBIOl,
input
CORETSE_AHBooI,
input
CORETSE_AHBlOl,
input
CORETSE_AHBoOl,
input
[
1
:
0
]
CORETSE_AHBiOl,
input
[
31
:
0
]
CORETSE_AHBOIl,
output
CORETSE_AHBIIl,
output
[
1
:
0
]
CORETSE_AHBlIl,
output
[
31
:
2
]
CORETSE_AHBoIl,
output
CORETSE_AHBiIl,
output
[
31
:
0
]
CORETSE_AHBOll,
input
CORETSE_AHBIll,
input
CORETSE_AHBlll,
input
[
1
:
0
]
CORETSE_AHBoll,
input
[
31
:
0
]
CORETSE_AHBill,
output
CORETSE_AHBO0l,
output
[
1
:
0
]
CORETSE_AHBI0l,
output
[
31
:
2
]
CORETSE_AHBl0l,
output
CORETSE_AHBo0l,
output
[
31
:
0
]
CORETSE_AHBi0l,
input
CORETSE_AHBO1l,
output
CORETSE_AHBI1l,
output
CORETSE_AHBl1l,
output
CORETSE_AHBo1l,
input
CORETSE_AHBOl0,
input
CORETSE_AHBIl0,
input
CORETSE_AHBlI0,
input
CORETSE_AHBoI0,
input
CORETSE_AHBiI0,
output
CORETSE_AHBll0,
output
CORETSE_AHBol0,
output
CORETSE_AHBil0,
output
CORETSE_AHBO00,
output
CORETSE_AHBI00,
output
CORETSE_AHBi1l,
output
CORETSE_AHBOol,
output
CORETSE_AHBIol,
output
[
TABITS
-
1
:
0
]
CORETSE_AHBlol,
output
[
39
:
0
]
CORETSE_AHBool,
output
[
TABITS
-
1
:
0
]
CORETSE_AHBiol,
input
[
39
:
0
]
CORETSE_AHBOil,
output
CORETSE_AHBIil,
output
CORETSE_AHBlil,
output
CORETSE_AHBoil,
output
[
RABITS
-
1
:
0
]
CORETSE_AHBiil,
output
[
35
:
0
]
CORETSE_AHBOO0,
output
[
RABITS
-
1
:
0
]
CORETSE_AHBIO0,
input
[
35
:
0
]
CORETSE_AHBlO0,
input
[
31
:
0
]
CORETSE_AHBl00,
output
[
31
:
0
]
CORETSE_AHBo00,
output
[
1
:
0
]
CORETSE_AHBO0,
output
CORETSE_AHBI0,
output
CORETSE_AHBoO0,
output
CORETSE_AHBl0,
output
CORETSE_AHBiO0,
output
CORETSE_AHBOI0,
output
CORETSE_AHBII0,
output
[
7
:
0
]
CORETSE_AHBi00
)
;
wire
[
31
:
0
]
CORETSE_AHBllIl
;
wire
CORETSE_AHBolIl
;
wire
[
31
:
0
]
CORETSE_AHBO0Il
;
wire
CORETSE_AHBI0Il
;
wire
CORETSE_AHBilIl
;
wire
[
1
:
0
]
CORETSE_AHBoo01
;
wire
CORETSE_AHBI11oI
;
wire
CORETSE_AHBl11oI
;
wire
[
31
:
0
]
CORETSE_AHBiIIl
;
wire
CORETSE_AHBOlIl
;
wire
CORETSE_AHBoIIl
;
wire
CORETSE_AHBo1llI
;
wire
[
7
:
0
]
CORETSE_AHBiOIlI
;
wire
[
7
:
0
]
CORETSE_AHBIl0lI
;
wire
CORETSE_AHBo1o1I
;
wire
[
7
:
0
]
CORETSE_AHBI1IOI
;
wire
[
7
:
0
]
CORETSE_AHBOii0
;
wire
CORETSE_AHBlO0OI
;
wire
CORETSE_AHBIO0OI
;
wire
CORETSE_AHBo11oI
;
wire
CORETSE_AHBi11oI
;
wire
CORETSE_AHBIo1II
;
wire
[
15
:
0
]
CORETSE_AHBOo1oI
;
wire
CORETSE_AHBIo1oI
;
wire
CORETSE_AHBIIO1I
;
wire
[
79
:
0
]
CORETSE_AHBi1I0I
;
wire
[
31
:
0
]
CORETSE_AHBIOo
;
wire
CORETSE_AHBlOo
;
wire
CORETSE_AHBoOo
;
wire
[
1
:
0
]
CORETSE_AHBiOo
;
wire
CORETSE_AHBiIo
;
wire
CORETSE_AHBIlo
;
wire
CORETSE_AHBIIo
;
wire
CORETSE_AHBOIo
;
wire
[
1
:
0
]
CORETSE_AHBlIo
;
wire
CORETSE_AHBoIo
;
wire
CORETSE_AHBloo
;
wire
CORETSE_AHBooo
;
wire
[
31
:
0
]
CORETSE_AHBioo
;
wire
CORETSE_AHBOio
;
wire
CORETSE_AHBIio
;
wire
[
1
:
0
]
CORETSE_AHBlio
;
wire
CORETSE_AHBoio
;
wire
[
7
:
0
]
CORETSE_AHBiio
;
wire
CORETSE_AHBOOi
;
wire
CORETSE_AHBIOi
;
wire
CORETSE_AHBlOi
;
wire
CORETSE_AHBiOi
;
wire
CORETSE_AHBOIi
;
wire
CORETSE_AHBIIi
;
wire
CORETSE_AHBoOi
;
wire
CORETSE_AHBlIi
;
wire
CORETSE_AHBoIi
;
wire
CORETSE_AHBolo
;
wire
CORETSE_AHBOOo1
;
wire
CORETSE_AHBilo
;
wire
CORETSE_AHBO0o
;
wire
CORETSE_AHBI0o
;
wire
CORETSE_AHBIoo
;
wire
[
7
:
0
]
CORETSE_AHBo0o
;
wire
CORETSE_AHBi0o
;
wire
CORETSE_AHBO1o
;
wire
CORETSE_AHBI1o
;
wire
CORETSE_AHBiOo1
;
wire
CORETSE_AHBo1o
;
wire
[
32
:
0
]
CORETSE_AHBl1o
;
wire
CORETSE_AHBIOo1
;
wire
[
51
:
0
]
CORETSE_AHBlOo1
;
wire
CORETSE_AHBIl00
;
wire
CORETSE_AHBi1o
;
wire
CORETSE_AHBOl00
;
wire
CORETSE_AHBiI00
;
wire
[
8
:
0
]
CORETSE_AHBIIo1
;
wire
CORETSE_AHBlIo1
;
wire
[
15
:
0
]
CORETSE_AHBOii1
;
wire
CORETSE_AHBIi1
;
wire
CORETSE_AHBli1
;
wire
[
7
:
0
]
CORETSE_AHBoi1
;
wire
[
31
:
0
]
CORETSE_AHBii1
;
wire
CORETSE_AHBI1i
;
wire
CORETSE_AHBlo1oI
;
wire
CORETSE_AHBoo1oI
;
wire
[
31
:
0
]
CORETSE_AHBO1i
;
wire
[
31
:
0
]
CORETSE_AHBio1oI
;
wire
[
31
:
0
]
CORETSE_AHBOi1oI
;
wire
[
31
:
0
]
CORETSE_AHBIi1oI
;
wire
CORETSE_AHBlOIi
;
wire
CORETSE_AHBoiOi
;
wire
CORETSE_AHBO1Ol
;
wire
CORETSE_AHBI1Ol
;
wire
[
31
:
0
]
CORETSE_AHBl1Ol
;
wire
CORETSE_AHBo1Ol
;
wire
CORETSE_AHBi1Ol
;
wire
[
1
:
0
]
CORETSE_AHBOoOl
;
wire
CORETSE_AHBli1oI
;
wire
CORETSE_AHBoi1oI
;
wire
[
47
:
0
]
CORETSE_AHBll00
;
wire
CORETSE_AHBol00
;
wire
CORETSE_AHBil00
;
wire
CORETSE_AHBI000
;
wire
CORETSE_AHBO000
;
wire
CORETSE_AHBii1oI
;
wire
CORETSE_AHBOOooI
;
wire
CORETSE_AHBOoOi
;
wire
[
5
:
0
]
CORETSE_AHBii0oI
;
wire
[
31
:
0
]
CORETSE_AHBOO1oI
;
wire
[
31
:
0
]
CORETSE_AHBIO1oI
;
wire
[
31
:
0
]
CORETSE_AHBlO1oI
;
wire
[
31
:
0
]
CORETSE_AHBoO1oI
;
wire
[
31
:
0
]
CORETSE_AHBii
,
CORETSE_AHBOOI
;
assign
CORETSE_AHBo00
=
CORETSE_AHBii
;
assign
CORETSE_AHBOOI
=
CORETSE_AHBl00
;
assign
CORETSE_AHBi1l
=
CORETSE_AHBloI
;
assign
CORETSE_AHBOol
=
CORETSE_AHBO0I
;
assign
CORETSE_AHBIil
=
CORETSE_AHBI0I
;
assign
CORETSE_AHBlil
=
CORETSE_AHBloI
;
assign
CORETSE_AHBO0
=
CORETSE_AHBoo01
;
generate
if
(
CORETSE_AHBiOI
==
0
)
begin
assign
CORETSE_AHBo1llI
=
1
'b
0
;
assign
CORETSE_AHBiOIlI
=
8
'b
0
;
assign
CORETSE_AHBIl0lI
=
8
'b
0
;
assign
CORETSE_AHBo1o1I
=
1
'b
0
;
assign
CORETSE_AHBI1IOI
=
8
'b
0
;
assign
CORETSE_AHBOii0
=
8
'b
0
;
assign
CORETSE_AHBlO0OI
=
1
'b
0
;
assign
CORETSE_AHBIO0OI
=
1
'b
0
;
assign
CORETSE_AHBo11oI
=
1
'b
0
;
assign
CORETSE_AHBi11oI
=
1
'b
0
;
assign
CORETSE_AHBIo1II
=
1
'b
0
;
assign
CORETSE_AHBOo1oI
=
8
'b
0
;
assign
CORETSE_AHBIo1oI
=
1
'b
0
;
assign
CORETSE_AHBIIO1I
=
1
'b
0
;
assign
CORETSE_AHBi1I0I
=
80
'b
0
;
end
endgenerate
mahbe_dual
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
,
.CORETSE_AHBOII
(
CORETSE_AHBOII
)
)
CORETSE_AHBIOooI
(
.CORETSE_AHBl1Il
(
CORETSE_AHBIoI
)
,
.HCLK
(
CORETSE_AHBloI
)
,
.CORETSE_AHBi0ll
(
CORETSE_AHBloo
)
,
.CORETSE_AHBO1ll
(
CORETSE_AHBooo
)
,
.CORETSE_AHBI1ll
(
CORETSE_AHBI1Ol
)
,
.CORETSE_AHBl1ll
(
CORETSE_AHBo1Ol
)
,
.CORETSE_AHBo1ll
(
CORETSE_AHBi1Ol
)
,
.CORETSE_AHBi1ll
(
CORETSE_AHBl1Ol
)
,
.CORETSE_AHBOoll
(
CORETSE_AHBOoOl
)
,
.CORETSE_AHBIiOl
(
CORETSE_AHBO1i
)
,
.CORETSE_AHBliOl
(
CORETSE_AHBI1i
)
,
.CORETSE_AHBO1l0
(
CORETSE_AHBlOIi
)
,
.CORETSE_AHBloI0
(
CORETSE_AHBioI
)
,
.CORETSE_AHBooI0
(
CORETSE_AHBOiI
)
,
.CORETSE_AHBioI0
(
CORETSE_AHBIiI
)
,
.CORETSE_AHBOiI0
(
CORETSE_AHBliI
)
,
.CORETSE_AHBIiI0
(
CORETSE_AHBoiI
)
,
.CORETSE_AHBliI0
(
CORETSE_AHBiiI
)
,
.CORETSE_AHBoiI0
(
CORETSE_AHBOOl
)
,
.CORETSE_AHBiiI0
(
CORETSE_AHBIOl
)
,
.CORETSE_AHBOOl0
(
CORETSE_AHBooI
)
,
.CORETSE_AHBIOl0
(
CORETSE_AHBlOl
)
,
.CORETSE_AHBoOl0
(
CORETSE_AHBiOl
)
,
.CORETSE_AHBiOl0
(
CORETSE_AHBOIl
)
,
.CORETSE_AHBOll0
(
CORETSE_AHBIll
)
,
.CORETSE_AHBlll0
(
CORETSE_AHBoll
)
,
.CORETSE_AHBoll0
(
CORETSE_AHBill
)
,
.CORETSE_AHBOIl0
(
CORETSE_AHBIIl
)
,
.CORETSE_AHBlOl0
(
CORETSE_AHBoOl
)
,
.CORETSE_AHBIIl0
(
CORETSE_AHBlIl
)
,
.CORETSE_AHBlIl0
(
CORETSE_AHBoIl
)
,
.CORETSE_AHBoIl0
(
CORETSE_AHBiIl
)
,
.CORETSE_AHBiIl0
(
CORETSE_AHBOll
)
,
.CORETSE_AHBill0
(
CORETSE_AHBO0l
)
,
.CORETSE_AHBIll0
(
CORETSE_AHBlll
)
,
.CORETSE_AHBO0l0
(
CORETSE_AHBI0l
)
,
.CORETSE_AHBI0l0
(
CORETSE_AHBl0l
)
,
.CORETSE_AHBl0l0
(
CORETSE_AHBo0l
)
,
.CORETSE_AHBo0l0
(
CORETSE_AHBi0l
)
,
.CORETSE_AHBiIll
(
CORETSE_AHBiIo
)
,
.CORETSE_AHBOlll
(
CORETSE_AHBlOo
)
,
.CORETSE_AHBIlll
(
CORETSE_AHBoOo
)
,
.CORETSE_AHBllll
(
CORETSE_AHBIOo
)
,
.CORETSE_AHBolll
(
CORETSE_AHBiOo
)
,
.CORETSE_AHBilll
(
CORETSE_AHBO1Ol
)
,
.CORETSE_AHBO0ll
(
CORETSE_AHBIIo
)
,
.CORETSE_AHBI0ll
(
CORETSE_AHBOIo
)
,
.CORETSE_AHBl0ll
(
CORETSE_AHBlIo
)
,
.CORETSE_AHBo0ll
(
CORETSE_AHBoIo
)
,
.CORETSE_AHBioOl
(
CORETSE_AHBIi1
)
,
.CORETSE_AHBIoll
(
CORETSE_AHBli1
)
,
.CORETSE_AHBOiOl
(
CORETSE_AHBoi1
)
,
.CORETSE_AHBloll
(
CORETSE_AHBii1
)
,
.CORETSE_AHBi0l0
(
CORETSE_AHBoiOi
)
,
.CORETSE_AHBI1l0
(
CORETSE_AHBii0oI
)
,
.CORETSE_AHBl1l0
(
CORETSE_AHBOO1oI
)
,
.CORETSE_AHBo1l0
(
CORETSE_AHBIO1oI
)
,
.CORETSE_AHBi1l0
(
CORETSE_AHBlO1oI
)
,
.CORETSE_AHBOol0
(
CORETSE_AHBoO1oI
)
,
.CORETSE_AHBl00
(
CORETSE_AHBOOI
)
,
.CORETSE_AHBo00
(
CORETSE_AHBii
)
,
.CORETSE_AHBIIll
(
CORETSE_AHBOii1
)
,
.CORETSE_AHBoIIl
(
CORETSE_AHBoIIl
)
,
.CORETSE_AHBiIIl
(
CORETSE_AHBiIIl
)
,
.CORETSE_AHBOlIl
(
CORETSE_AHBOlIl
)
,
.CORETSE_AHBIlIl
(
CORETSE_AHBIlIl
)
,
.CORETSE_AHBllIl
(
CORETSE_AHBllIl
)
,
.CORETSE_AHBolIl
(
CORETSE_AHBolIl
)
,
.CORETSE_AHBilIl
(
CORETSE_AHBilIl
)
,
.CORETSE_AHBO0Il
(
CORETSE_AHBO0Il
)
,
.CORETSE_AHBI0Il
(
CORETSE_AHBI0Il
)
,
.CORETSE_AHBooll
(
CORETSE_AHBoi1oI
)
)
;
arfque
CORETSE_AHBlOooI
(
.CORETSE_AHBo0Ol
(
CORETSE_AHBloI
)
,
.CORETSE_AHBi0Ol
(
CORETSE_AHBIoI
)
,
.CORETSE_AHBoio
(
CORETSE_AHBoio
)
,
.CORETSE_AHBioo
(
CORETSE_AHBioo
)
,
.CORETSE_AHBOio
(
CORETSE_AHBOio
)
,
.CORETSE_AHBIio
(
CORETSE_AHBIio
)
,
.CORETSE_AHBlio
(
CORETSE_AHBlio
)
,
.CORETSE_AHBO1Ol
(
CORETSE_AHBO1Ol
)
,
.CORETSE_AHBIlo
(
CORETSE_AHBIlo
)
,
.CORETSE_AHBI1Ol
(
CORETSE_AHBI1Ol
)
,
.CORETSE_AHBl1Ol
(
CORETSE_AHBl1Ol
)
,
.CORETSE_AHBo1Ol
(
CORETSE_AHBo1Ol
)
,
.CORETSE_AHBi1Ol
(
CORETSE_AHBi1Ol
)
,
.CORETSE_AHBOoOl
(
CORETSE_AHBOoOl
)
)
;
assign
CORETSE_AHBi1o
=
(
!
CORETSE_AHBIl00
&
!
CORETSE_AHBOl00
&
!
CORETSE_AHBiI00
)
;
amcxfif
#
(
.TABITS
(
TABITS
)
,
.RABITS
(
RABITS
)
,
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
)
CORETSE_AHBoOooI
(
.CORETSE_AHBIi0
(
~
CORETSE_AHBIoI
)
,
.CORETSE_AHBoo1
(
CORETSE_AHBl0I
)
,
.CORETSE_AHBio1
(
~
CORETSE_AHBIoI
)
,
.CORETSE_AHBOi1
(
CORETSE_AHBloI
)
,
.CORETSE_AHBIi1
(
CORETSE_AHBIi1
)
,
.CORETSE_AHBli1
(
CORETSE_AHBli1
)
,
.CORETSE_AHBoi1
(
CORETSE_AHBoi1
)
,
.CORETSE_AHBii1
(
CORETSE_AHBii1
)
,
.CORETSE_AHBOOo
(
CORETSE_AHBloI
)
,
.CORETSE_AHBIOo
(
CORETSE_AHBIOo
)
,
.CORETSE_AHBlOo
(
CORETSE_AHBlOo
)
,
.CORETSE_AHBoOo
(
CORETSE_AHBoOo
)
,
.CORETSE_AHBiOo
(
CORETSE_AHBiOo
)
,
.CORETSE_AHBOIo
(
CORETSE_AHBOIo
)
,
.CORETSE_AHBIIo
(
CORETSE_AHBIIo
)
,
.CORETSE_AHBlIo
(
CORETSE_AHBlIo
)
,
.CORETSE_AHBoIo
(
CORETSE_AHBoIo
)
,
.CORETSE_AHBiIo
(
CORETSE_AHBiIo
)
,
.CORETSE_AHBOlo
(
CORETSE_AHBloI
)
,
.CORETSE_AHBIlo
(
CORETSE_AHBIlo
)
,
.CORETSE_AHBoi0
(
CORETSE_AHBO0I
)
,
.CORETSE_AHBllo
(
1
'b
1
)
,
.CORETSE_AHBolo
(
CORETSE_AHBolo
)
,
.CORETSE_AHBilo
(
CORETSE_AHBilo
)
,
.CORETSE_AHBO0o
(
CORETSE_AHBO0o
)
,
.CORETSE_AHBI0o
(
CORETSE_AHBI0o
)
,
.CORETSE_AHBii0
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBl0o
(
1
'b
1
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBo0o
)
,
.CORETSE_AHBi0o
(
CORETSE_AHBi0o
)
,
.CORETSE_AHBO1o
(
CORETSE_AHBO1o
)
,
.CORETSE_AHBI1o
(
CORETSE_AHBI1o
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBi1o
(
CORETSE_AHBi1o
)
,
.CORETSE_AHBOoo
(
CORETSE_AHBOOooI
)
,
.CORETSE_AHBIoo
(
CORETSE_AHBIoo
)
,
.CORETSE_AHBloo
(
CORETSE_AHBloo
)
,
.CORETSE_AHBooo
(
CORETSE_AHBooo
)
,
.CORETSE_AHBioo
(
CORETSE_AHBioo
)
,
.CORETSE_AHBOio
(
CORETSE_AHBOio
)
,
.CORETSE_AHBIio
(
CORETSE_AHBIio
)
,
.CORETSE_AHBlio
(
CORETSE_AHBlio
)
,
.CORETSE_AHBoio
(
CORETSE_AHBoio
)
,
.CORETSE_AHBiio
(
CORETSE_AHBiio
)
,
.CORETSE_AHBOOi
(
CORETSE_AHBOOi
)
,
.CORETSE_AHBIOi
(
CORETSE_AHBIOi
)
,
.CORETSE_AHBlOi
(
CORETSE_AHBlOi
)
,
.CORETSE_AHBoOi
(
CORETSE_AHBoOi
)
,
.CORETSE_AHBiOi
(
CORETSE_AHBiOi
)
,
.CORETSE_AHBOIi
(
CORETSE_AHBOIi
)
,
.CORETSE_AHBIIi
(
CORETSE_AHBIIi
)
,
.CORETSE_AHBlIi
(
CORETSE_AHBlIi
)
,
.CORETSE_AHBoIi
(
CORETSE_AHBoIi
)
,
.CORETSE_AHBiIi
(
CORETSE_AHBiIi
)
,
.CORETSE_AHBOli
(
CORETSE_AHBIol
)
,
.CORETSE_AHBIli
(
CORETSE_AHBlol
)
,
.CORETSE_AHBlli
(
CORETSE_AHBool
)
,
.CORETSE_AHBoli
(
CORETSE_AHBiol
)
,
.CORETSE_AHBili
(
CORETSE_AHBOil
)
,
.CORETSE_AHBO0i
(
CORETSE_AHBoil
)
,
.CORETSE_AHBI0i
(
CORETSE_AHBiil
)
,
.CORETSE_AHBl0i
(
CORETSE_AHBOO0
)
,
.CORETSE_AHBo0i
(
CORETSE_AHBIO0
)
,
.CORETSE_AHBi0i
(
CORETSE_AHBlO0
)
,
.CORETSE_AHBO1i
(
CORETSE_AHBio1oI
)
,
.CORETSE_AHBI1i
(
CORETSE_AHBlo1oI
)
)
;
pe_mcxmac
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
,
.CORETSE_AHBiOI
(
CORETSE_AHBiOI
)
)
CORETSE_AHBiOooI
(
.CORETSE_AHBO111
(
1
'b
0
)
,
.CORETSE_AHBI111
(
1
'b
0
)
,
.CORETSE_AHBl111
(
1
'b
0
)
,
.CORETSE_AHBiOO1
(
1
'b
0
)
,
.CORETSE_AHBoi0
(
CORETSE_AHBO0I
)
,
.CORETSE_AHBllo
(
1
'b
1
)
,
.CORETSE_AHBo111
(
1
'b
0
)
,
.CORETSE_AHBii0
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBl0o
(
1
'b
1
)
,
.CORETSE_AHBol
(
CORETSE_AHBo0I
)
,
.CORETSE_AHBll
(
CORETSE_AHBi0I
)
,
.CORETSE_AHBo01
(
CORETSE_AHBO1l
)
,
.CORETSE_AHBiio
(
CORETSE_AHBiio
)
,
.CORETSE_AHBiOi
(
CORETSE_AHBiOi
)
,
.CORETSE_AHBOIi
(
CORETSE_AHBOIi
)
,
.CORETSE_AHBIIi
(
CORETSE_AHBIIi
)
,
.CORETSE_AHBoOi
(
CORETSE_AHBoOi
)
,
.CORETSE_AHBlIi
(
CORETSE_AHBlIi
)
,
.CORETSE_AHBi111
(
{
16
{
CORETSE_AHBoIi
}
}
)
,
.CORETSE_AHBiIi
(
CORETSE_AHBiIi
)
,
.CORETSE_AHBI000
(
CORETSE_AHBI000
)
,
.CORETSE_AHBol00
(
CORETSE_AHBol00
)
,
.CORETSE_AHBil00
(
CORETSE_AHBil00
)
,
.CORETSE_AHBO000
(
CORETSE_AHBO000
)
,
.CORETSE_AHBOo11
(
CORETSE_AHBOo11
)
,
.CORETSE_AHBIo11
(
CORETSE_AHBIo11
)
,
.CORETSE_AHBoo01
(
CORETSE_AHBoo01
)
,
.CORETSE_AHBlo11
(
CORETSE_AHBlo11
)
,
.CORETSE_AHBiI
(
CORETSE_AHBO1I
)
,
.CORETSE_AHBlI
(
CORETSE_AHBI1I
)
,
.CORETSE_AHBIl
(
CORETSE_AHBl1I
)
,
.CORETSE_AHBlOi
(
CORETSE_AHBlOi
)
,
.CORETSE_AHBOOi
(
CORETSE_AHBOOi
)
,
.CORETSE_AHBoo11
(
1
'b
0
)
,
.CORETSE_AHBIOi
(
CORETSE_AHBIOi
)
,
.CORETSE_AHBio1
(
~
CORETSE_AHBIoI
)
,
.CORETSE_AHBOi1
(
CORETSE_AHBloI
)
,
.CORETSE_AHBIi1
(
CORETSE_AHBIi1
)
,
.CORETSE_AHBli1
(
CORETSE_AHBli1
)
,
.CORETSE_AHBoi1
(
CORETSE_AHBoi1
)
,
.CORETSE_AHBii1
(
CORETSE_AHBii1
)
,
.CORETSE_AHBoo1
(
CORETSE_AHBl0I
)
,
.CORETSE_AHBll00
(
CORETSE_AHBll00
)
,
.CORETSE_AHBio11
(
CORETSE_AHBloI
)
,
.CORETSE_AHBOi11
(
5
'b
0
)
,
.CORETSE_AHBIi11
(
)
,
.CORETSE_AHBli11
(
)
,
.CORETSE_AHBoi11
(
)
,
.CORETSE_AHBii11
(
)
,
.CORETSE_AHBoI
(
CORETSE_AHBo1I
)
,
.CORETSE_AHBII
(
CORETSE_AHBi1I
)
,
.CORETSE_AHBOl
(
CORETSE_AHBOoI
)
,
.CORETSE_AHBi01
(
CORETSE_AHBI1l
)
,
.CORETSE_AHBO11
(
CORETSE_AHBl1l
)
,
.CORETSE_AHBI11
(
CORETSE_AHBo1l
)
,
.CORETSE_AHBolo
(
CORETSE_AHBolo
)
,
.CORETSE_AHBOOo1
(
CORETSE_AHBOOo1
)
,
.CORETSE_AHBO0o
(
CORETSE_AHBO0o
)
,
.CORETSE_AHBilo
(
CORETSE_AHBilo
)
,
.CORETSE_AHBI0o
(
CORETSE_AHBI0o
)
,
.CORETSE_AHBIOo1
(
CORETSE_AHBIOo1
)
,
.CORETSE_AHBlOo1
(
CORETSE_AHBlOo1
)
,
.CORETSE_AHBoOo1
(
CORETSE_AHBOIooI
)
,
.CORETSE_AHBIoo
(
CORETSE_AHBIoo
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBo0o
)
,
.CORETSE_AHBi0o
(
CORETSE_AHBi0o
)
,
.CORETSE_AHBO1o
(
CORETSE_AHBO1o
)
,
.CORETSE_AHBI1o
(
CORETSE_AHBI1o
)
,
.CORETSE_AHBiOo1
(
CORETSE_AHBiOo1
)
,
.CORETSE_AHBOIo1
(
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
)
,
.CORETSE_AHBIIo1
(
CORETSE_AHBIIo1
)
,
.CORETSE_AHBlIo1
(
CORETSE_AHBlIo1
)
,
.CORETSE_AHBiI00
(
CORETSE_AHBiI00
)
,
.CORETSE_AHBOl00
(
CORETSE_AHBOl00
)
,
.CORETSE_AHBIl00
(
CORETSE_AHBIl00
)
,
.CORETSE_AHBO1i
(
CORETSE_AHBOi1oI
)
,
.CORETSE_AHBI1i
(
CORETSE_AHBoo1oI
)
,
.CORETSE_AHBoIo1
(
CORETSE_AHBI0
)
,
.CORETSE_AHBiIo1
(
CORETSE_AHBoO0
)
,
.CORETSE_AHBOlo1
(
CORETSE_AHBl0
)
,
.CORETSE_AHBIlo1
(
CORETSE_AHBiO0
)
,
.CORETSE_AHBO0o1
(
CORETSE_AHBOii1
)
,
.CORETSE_AHBI0o1
(
CORETSE_AHBo1llI
)
,
.CORETSE_AHBl0o1
(
CORETSE_AHBiOIlI
)
,
.CORETSE_AHBo0o1
(
CORETSE_AHBIl0lI
)
,
.CORETSE_AHBi0o1
(
CORETSE_AHBo1o1I
)
,
.CORETSE_AHBO1o1
(
CORETSE_AHBI1IOI
)
,
.CORETSE_AHBI1o1
(
CORETSE_AHBOii0
)
,
.CORETSE_AHBl1o1
(
CORETSE_AHBlO0OI
)
,
.CORETSE_AHBo1o1
(
CORETSE_AHBIO0OI
)
,
.CORETSE_AHBi1o1
(
CORETSE_AHBo11oI
)
,
.CORETSE_AHBOoo1
(
CORETSE_AHBi11oI
)
,
.CORETSE_AHBIoo1
(
CORETSE_AHBIo1II
)
,
.CORETSE_AHBloo1
(
CORETSE_AHBOo1oI
)
,
.CORETSE_AHBooo1
(
CORETSE_AHBIo1oI
)
,
.CORETSE_AHBOio1
(
CORETSE_AHBIIO1I
)
,
.CORETSE_AHBioo1
(
CORETSE_AHBi1I0I
)
,
.CORETSE_AHBllo1
(
)
,
.CORETSE_AHBolo1
(
CORETSE_AHBOI0
)
,
.CORETSE_AHBilo1
(
CORETSE_AHBII0
)
,
.CORETSE_AHBIio1
(
CORETSE_AHBIio1
)
,
.CORETSE_AHBlio1
(
CORETSE_AHBlio1
)
,
.CORETSE_AHBoio1
(
)
,
.CORETSE_AHBiio1
(
)
)
;
generate
if
(
CORETSE_AHBiOI
==
1
)
begin
:
CORETSE_AHBIIooI
ptp_top
#
(
.CORETSE_AHBIII
(
CORETSE_AHBIII
)
,
.CORETSE_AHBlII
(
CORETSE_AHBlII
)
,
.CORETSE_AHBoII
(
CORETSE_AHBoII
)
,
.CORETSE_AHBiII
(
CORETSE_AHBiII
)
,
.CORETSE_AHBOlI
(
CORETSE_AHBOlI
)
,
.CORETSE_AHBIlI
(
CORETSE_AHBIlI
)
,
.CORETSE_AHBllI
(
CORETSE_AHBllI
)
,
.CORETSE_AHBolI
(
CORETSE_AHBolI
)
)
CORETSE_AHBlIooI
(
.CORETSE_AHBiil0
(
CORETSE_AHBloI
)
,
.CORETSE_AHBi10lI
(
~
CORETSE_AHBIoI
)
,
.CORETSE_AHBOl0
(
CORETSE_AHBOl0
)
,
.CORETSE_AHBOo0lI
(
~
CORETSE_AHBIoI
)
,
.CORETSE_AHBl0I
(
CORETSE_AHBl0I
)
,
.CORETSE_AHBIl0
(
CORETSE_AHBIl0
)
,
.CORETSE_AHBOI01I
(
CORETSE_AHBO0I
)
,
.CORETSE_AHBII01I
(
CORETSE_AHBIio1
)
,
.CORETSE_AHBlI01I
(
1
'b
1
)
,
.CORETSE_AHBoI01I
(
CORETSE_AHBo1llI
)
,
.CORETSE_AHBoIo0I
(
CORETSE_AHBoo01
)
,
.CORETSE_AHBiI01I
(
CORETSE_AHBiOIlI
)
,
.CORETSE_AHBOl01I
(
CORETSE_AHBIl0lI
)
,
.CORETSE_AHBi1O1I
(
CORETSE_AHBo1o1I
)
,
.CORETSE_AHBOOo0I
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBiOo0I
(
1
'b
1
)
,
.CORETSE_AHBIOo0I
(
CORETSE_AHBlio1
)
,
.CORETSE_AHBlo0lI
(
CORETSE_AHBoIIl
)
,
.CORETSE_AHBoo0lI
(
CORETSE_AHBli1
)
,
.CORETSE_AHBoO00
(
CORETSE_AHBoi1
[
4
:
0
]
)
,
.CORETSE_AHBioo1I
(
CORETSE_AHBii1
)
,
.CORETSE_AHBOIo0I
(
CORETSE_AHBOii0
)
,
.CORETSE_AHBIIo0I
(
CORETSE_AHBI1IOI
)
,
.CORETSE_AHBOoO1I
(
CORETSE_AHBlO0OI
)
,
.CORETSE_AHBlIo0I
(
CORETSE_AHBIO0OI
)
,
.CORETSE_AHBiIo0I
(
CORETSE_AHBo11oI
)
,
.CORETSE_AHBlI0
(
CORETSE_AHBlI0
)
,
.CORETSE_AHBoI0
(
CORETSE_AHBoI0
)
,
.CORETSE_AHBiI0
(
CORETSE_AHBiI0
)
,
.CORETSE_AHBOio1I
(
CORETSE_AHBiIIl
)
,
.CORETSE_AHBIio1I
(
)
,
.CORETSE_AHBOl1lI
(
CORETSE_AHBl11oI
)
,
.CORETSE_AHBlio1I
(
CORETSE_AHBOlIl
)
,
.CORETSE_AHBO001I
(
CORETSE_AHBi11oI
)
,
.CORETSE_AHBl001I
(
CORETSE_AHBIo1II
)
,
.CORETSE_AHBo001I
(
CORETSE_AHBOo1oI
)
,
.CORETSE_AHBI101I
(
CORETSE_AHBIo1oI
)
,
.CORETSE_AHBO101I
(
CORETSE_AHBIIO1I
)
,
.CORETSE_AHBoio1I
(
CORETSE_AHBi1I0I
)
,
.CORETSE_AHBll0
(
CORETSE_AHBll0
)
,
.CORETSE_AHBol0
(
CORETSE_AHBol0
)
,
.CORETSE_AHBil0
(
CORETSE_AHBil0
)
,
.CORETSE_AHBO00
(
CORETSE_AHBO00
)
,
.CORETSE_AHBI00
(
CORETSE_AHBI00
)
)
;
end
else
begin
assign
CORETSE_AHBl11oI
=
1
'b
0
;
assign
CORETSE_AHBiIIl
=
32
'b
0
;
assign
CORETSE_AHBOlIl
=
1
'b
0
;
end
endgenerate
assign
CORETSE_AHBI11oI
=
1
'b
0
;
assign
CORETSE_AHBllIl
=
32
'b
0
;
assign
CORETSE_AHBolIl
=
1
'b
0
;
assign
CORETSE_AHBO0Il
=
32
'b
0
;
assign
CORETSE_AHBI0Il
=
1
'b
0
;
assign
CORETSE_AHBoIooI
=
1
'b
0
;
assign
CORETSE_AHBiIooI
=
1
'b
0
;
generate
if
(
MCXMAC_STATS_ON
==
1
)
begin
:
CORETSE_AHBOlooI
wire
CORETSE_AHBo1Oi
,
CORETSE_AHBi1Oi
,
CORETSE_AHBIlooI
,
CORETSE_AHBllooI
;
assign
CORETSE_AHBo1Oi
=
CORETSE_AHBloI
;
assign
CORETSE_AHBi1Oi
=
~
CORETSE_AHBIoI
;
sib_sync_pulse
CORETSE_AHBolooI
(
.CORETSE_AHBO0I
(
CORETSE_AHBO0I
)
,
.CORETSE_AHBooloI
(
!
CORETSE_AHBIio1
)
,
.CORETSE_AHBioloI
(
CORETSE_AHBIOo1
)
,
.CORETSE_AHBI0I
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBOiloI
(
~
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBIiloI
(
CORETSE_AHBIlooI
)
,
.CORETSE_AHBliloI
(
)
)
;
sib_sync_pulse
CORETSE_AHBilooI
(
.CORETSE_AHBO0I
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBooloI
(
!
CORETSE_AHBlio1
)
,
.CORETSE_AHBioloI
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBI0I
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBOiloI
(
~
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBIiloI
(
CORETSE_AHBllooI
)
,
.CORETSE_AHBliloI
(
)
)
;
pemstat
CORETSE_AHBO0ooI
(
.CORETSE_AHBo1Oi
(
CORETSE_AHBo1Oi
)
,
.CORETSE_AHBi1Oi
(
CORETSE_AHBi1Oi
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
[
30
:
0
]
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBllooI
)
,
.CORETSE_AHBlOo1
(
CORETSE_AHBlOo1
)
,
.CORETSE_AHBIOo1
(
CORETSE_AHBIlooI
)
,
.CORETSE_AHBOoOi
(
CORETSE_AHBOoOi
)
,
.CORETSE_AHBIoOi
(
1
'b
0
)
,
.CORETSE_AHBloOi
(
1
'b
0
)
,
.CORETSE_AHBooOi
(
CORETSE_AHBOo11
)
,
.CORETSE_AHBioOi
(
CORETSE_AHBIo11
)
,
.CORETSE_AHBOiOi
(
CORETSE_AHBlo11
)
,
.CORETSE_AHBIiOi
(
1
'b
0
)
,
.CORETSE_AHBliOi
(
CORETSE_AHBoi1
[
6
:
0
]
)
,
.CORETSE_AHBoiOi
(
CORETSE_AHBoiOi
)
,
.CORETSE_AHBiiOi
(
CORETSE_AHBli1
)
,
.CORETSE_AHBOOIi
(
CORETSE_AHBii1
)
,
.CORETSE_AHBIOIi
(
CORETSE_AHBIi1oI
)
,
.CORETSE_AHBlOIi
(
CORETSE_AHBlOIi
)
,
.CORETSE_AHBoOIi
(
CORETSE_AHBli1oI
)
)
;
end
else
begin
assign
CORETSE_AHBIi1oI
=
32
'b
0
;
assign
CORETSE_AHBlOIi
=
1
'b
0
;
assign
CORETSE_AHBli1oI
=
1
'b
0
;
end
endgenerate
assign
CORETSE_AHBO1i
=
CORETSE_AHBOi1oI
|
CORETSE_AHBio1oI
|
CORETSE_AHBIi1oI
;
assign
CORETSE_AHBI1i
=
CORETSE_AHBoo1oI
|
CORETSE_AHBlo1oI
|
CORETSE_AHBlOIi
;
assign
CORETSE_AHBi00
=
{
3
'b
0
,
CORETSE_AHBI11oI
,
CORETSE_AHBii1oI
,
CORETSE_AHBl11oI
,
CORETSE_AHBli1oI
,
CORETSE_AHBoi1oI
}
;
generate
if
(
MCXMAC_WOL_ON
==
1
)
begin
:
CORETSE_AHBI0ooI
assign
CORETSE_AHBii1oI
=
CORETSE_AHBI000
&
CORETSE_AHBil00
;
mmcxwol
CORETSE_AHBl0ooI
(
.CORETSE_AHBii0
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBl0o
(
1
'b
1
)
,
.CORETSE_AHBl0II
(
CORETSE_AHBlio1
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBo0o
)
,
.CORETSE_AHBi0o
(
CORETSE_AHBi0o
)
,
.CORETSE_AHBO1o
(
CORETSE_AHBO1o
)
,
.CORETSE_AHBI1o
(
CORETSE_AHBI1o
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
[
22
:
20
]
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBiI00
(
CORETSE_AHBiI00
)
,
.CORETSE_AHBOl00
(
CORETSE_AHBOl00
)
,
.CORETSE_AHBIl00
(
CORETSE_AHBIl00
)
,
.CORETSE_AHBll00
(
CORETSE_AHBll00
)
,
.CORETSE_AHBol00
(
CORETSE_AHBol00
)
,
.CORETSE_AHBil00
(
CORETSE_AHBil00
)
,
.CORETSE_AHBO000
(
CORETSE_AHBO000
)
,
.CORETSE_AHBI000
(
CORETSE_AHBI000
)
)
;
end
else
begin
assign
CORETSE_AHBI000
=
1
'b
0
;
assign
CORETSE_AHBii1oI
=
1
'b
0
;
end
endgenerate
generate
if
(
MCXMAC_SAL_ON
==
1
)
begin
:
CORETSE_AHBo0ooI
si_sal
CORETSE_AHBi0ooI
(
.CORETSE_AHBioOoI
(
CORETSE_AHBI0I
)
,
.CORETSE_AHBOiOoI
(
!
CORETSE_AHBlio1
)
,
.CORETSE_AHBIiOoI
(
CORETSE_AHBIIo1
[
8
:
2
]
)
,
.CORETSE_AHBliOoI
(
CORETSE_AHBlIo1
)
,
.CORETSE_AHBoiOoI
(
CORETSE_AHBIl00
)
,
.CORETSE_AHBiiOoI
(
CORETSE_AHBOl00
)
,
.CORETSE_AHBOOIoI
(
CORETSE_AHBiI00
)
,
.CORETSE_AHBIOIoI
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBlOIoI
(
CORETSE_AHBii0oI
)
,
.CORETSE_AHBoOIoI
(
CORETSE_AHBOO1oI
)
,
.CORETSE_AHBiOIoI
(
CORETSE_AHBIO1oI
)
,
.CORETSE_AHBOIIoI
(
CORETSE_AHBlO1oI
)
,
.CORETSE_AHBIIIoI
(
CORETSE_AHBoO1oI
)
,
.CORETSE_AHBlIIoI
(
CORETSE_AHBOoOi
)
,
.CORETSE_AHBoIIoI
(
CORETSE_AHBOOooI
)
)
;
end
else
begin
assign
CORETSE_AHBOOooI
=
1
'b
0
;
assign
CORETSE_AHBOoOi
=
1
'b
0
;
end
endgenerate
endmodule
