// REVISION    : $Revision: 1.7 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxfif_hst
#
(
parameter
TABITS
=
12
,
parameter
RABITS
=
12
,
parameter
CORETSE_AHBIo1
=
32
,
parameter
CORETSE_AHBlo1
=
$clog2
(
CORETSE_AHBIo1
/
8
)
)
(
CORETSE_AHBio1
,
CORETSE_AHBOi1
,
CORETSE_AHBIi1
,
CORETSE_AHBli1
,
CORETSE_AHBoi1
,
CORETSE_AHBii1
,
CORETSE_AHBoOOI
,
CORETSE_AHBiOOI
,
CORETSE_AHBOIOI
,
CORETSE_AHBIIOI
,
CORETSE_AHBlIOI
,
CORETSE_AHBoIOI
,
CORETSE_AHBiIOI
,
CORETSE_AHBOlOI
,
CORETSE_AHBIlOI
,
CORETSE_AHBllOI
,
CORETSE_AHBolOI
,
CORETSE_AHBilOI
,
CORETSE_AHBO0OI
,
CORETSE_AHBI0OI
,
CORETSE_AHBl1OI
,
CORETSE_AHBo1OI
,
CORETSE_AHBi1OI
,
CORETSE_AHBl0OI
,
CORETSE_AHBo0OI
,
CORETSE_AHBi0OI
,
CORETSE_AHBO1OI
,
CORETSE_AHBI1OI
,
CORETSE_AHBOoOI
,
CORETSE_AHBIoOI
,
CORETSE_AHBloOI
,
CORETSE_AHBooOI
,
CORETSE_AHBioOI
,
CORETSE_AHBOiOI
,
CORETSE_AHBIiOI
,
CORETSE_AHBliOI
,
CORETSE_AHBoiOI
,
CORETSE_AHBiiOI
,
CORETSE_AHBOOII
,
CORETSE_AHBIOII
,
CORETSE_AHBlOII
,
CORETSE_AHBoOII
,
CORETSE_AHBiOII
,
CORETSE_AHBOIII
,
CORETSE_AHBIIII
,
CORETSE_AHBlIII
,
CORETSE_AHBoIII
,
CORETSE_AHBiIII
,
CORETSE_AHBOlII
,
CORETSE_AHBIlII
,
CORETSE_AHBllII
,
CORETSE_AHBolII
,
CORETSE_AHBO1i
,
CORETSE_AHBI1i
)
;
input
CORETSE_AHBio1
;
input
CORETSE_AHBOi1
;
input
CORETSE_AHBIi1
;
input
CORETSE_AHBli1
;
input
[
7
:
0
]
CORETSE_AHBoi1
;
input
[
31
:
0
]
CORETSE_AHBii1
;
input
CORETSE_AHBoOOI
;
input
CORETSE_AHBiOOI
;
input
CORETSE_AHBOIOI
;
input
CORETSE_AHBIIOI
;
input
CORETSE_AHBlIOI
;
input
CORETSE_AHBoIOI
;
input
CORETSE_AHBiIOI
;
input
[
TABITS
:
0
]
CORETSE_AHBOlOI
;
input
CORETSE_AHBIlOI
;
input
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBllOI
;
input
CORETSE_AHBolOI
;
input
[
RABITS
:
0
]
CORETSE_AHBilOI
;
input
CORETSE_AHBO0OI
;
input
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBI0OI
;
output
[
TABITS
:
0
]
CORETSE_AHBl1OI
;
output
[
TABITS
:
0
]
CORETSE_AHBo1OI
;
output
[
RABITS
-
1
:
0
]
CORETSE_AHBi1OI
;
output
[
15
:
0
]
CORETSE_AHBl0OI
;
output
[
RABITS
:
0
]
CORETSE_AHBo0OI
;
output
[
RABITS
:
0
]
CORETSE_AHBi0OI
;
output
CORETSE_AHBO1OI
;
output
CORETSE_AHBI1OI
;
output
[
17
:
0
]
CORETSE_AHBOoOI
;
output
[
17
:
0
]
CORETSE_AHBIoOI
;
output
CORETSE_AHBloOI
;
output
CORETSE_AHBooOI
;
output
CORETSE_AHBioOI
;
output
CORETSE_AHBOiOI
;
output
CORETSE_AHBIiOI
;
output
CORETSE_AHBliOI
;
output
CORETSE_AHBoiOI
;
output
CORETSE_AHBiiOI
;
output
CORETSE_AHBOOII
;
output
CORETSE_AHBIOII
;
output
CORETSE_AHBlOII
;
output
CORETSE_AHBoOII
;
output
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBiOII
;
output
CORETSE_AHBOIII
;
output
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIIII
;
output
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBlIII
;
output
CORETSE_AHBoIII
;
output
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBiIII
;
output
CORETSE_AHBOlII
;
output
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIlII
;
output
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBllII
;
output
CORETSE_AHBolII
;
output
[
31
:
0
]
CORETSE_AHBO1i
;
output
CORETSE_AHBI1i
;
reg
[
TABITS
:
0
]
CORETSE_AHBl1OI
;
reg
[
TABITS
:
0
]
CORETSE_AHBo1OI
;
reg
[
RABITS
-
1
:
0
]
CORETSE_AHBi1OI
;
reg
[
15
:
0
]
CORETSE_AHBl0OI
;
reg
[
RABITS
:
0
]
CORETSE_AHBo0OI
;
reg
[
RABITS
:
0
]
CORETSE_AHBi0OI
;
reg
CORETSE_AHBO1OI
;
reg
CORETSE_AHBI1OI
;
reg
[
17
:
0
]
CORETSE_AHBOoOI
;
reg
[
17
:
0
]
CORETSE_AHBIoOI
;
reg
CORETSE_AHBloOI
;
reg
CORETSE_AHBooOI
;
reg
CORETSE_AHBioOI
;
reg
CORETSE_AHBOiOI
;
reg
CORETSE_AHBIiOI
;
reg
CORETSE_AHBliOI
;
reg
CORETSE_AHBoiOI
;
reg
CORETSE_AHBiiOI
;
reg
CORETSE_AHBOOII
;
reg
CORETSE_AHBIOII
;
reg
CORETSE_AHBlOII
;
reg
CORETSE_AHBoOII
;
reg
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBiOII
;
reg
CORETSE_AHBOIII
;
reg
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIIII
;
reg
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBlIII
;
reg
CORETSE_AHBoIII
;
reg
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBiIII
;
reg
CORETSE_AHBOlII
;
reg
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIlII
;
reg
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBllII
;
reg
CORETSE_AHBolII
;
wire
[
31
:
0
]
CORETSE_AHBO1i
;
wire
CORETSE_AHBI1i
;
parameter
CORETSE_AHBIoII
=
1
;
parameter
CORETSE_AHBlOlI
=
{
(
TABITS
+
2
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBoOlI
=
{
(
15
-
TABITS
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBiOlI
=
{
(
30
-
TABITS
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBOIlI
=
{
(
TABITS
+
1
)
{
1
'b
1
}
}
;
parameter
CORETSE_AHBIIlI
=
{
(
RABITS
)
{
1
'b
1
}
}
;
parameter
CORETSE_AHBlIlI
=
{
(
RABITS
+
2
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBoIlI
=
{
(
16
-
RABITS
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBiIlI
=
{
(
15
-
RABITS
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBOllI
=
{
(
30
-
RABITS
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBIllI
=
{
(
RABITS
+
1
)
{
1
'b
1
}
}
;
parameter
CORETSE_AHBlllI
=
{
(
RABITS
+
1
)
{
1
'b
1
}
}
;
parameter
CORETSE_AHBollI
=
{
(
TABITS
+
1
)
{
1
'b
1
}
}
;
wire
CORETSE_AHBillI
;
wire
CORETSE_AHBO0lI
;
wire
CORETSE_AHBI0lI
;
wire
CORETSE_AHBl0lI
;
wire
CORETSE_AHBo0lI
;
wire
CORETSE_AHBi0lI
;
wire
CORETSE_AHBO1lI
;
wire
CORETSE_AHBI1lI
;
wire
CORETSE_AHBl1lI
;
wire
CORETSE_AHBo1lI
;
wire
CORETSE_AHBi1lI
;
wire
CORETSE_AHBOolI
;
wire
CORETSE_AHBIolI
;
wire
CORETSE_AHBlolI
;
wire
CORETSE_AHBoolI
;
wire
CORETSE_AHBiolI
;
wire
CORETSE_AHBOilI
;
wire
CORETSE_AHBIilI
;
wire
CORETSE_AHBlilI
;
wire
CORETSE_AHBoilI
;
wire
CORETSE_AHBiilI
;
wire
CORETSE_AHBOO0I
;
wire
CORETSE_AHBIO0I
;
wire
CORETSE_AHBlO0I
;
wire
CORETSE_AHBoO0I
;
wire
CORETSE_AHBiO0I
;
wire
CORETSE_AHBOI0I
;
wire
CORETSE_AHBII0I
;
wire
CORETSE_AHBlI0I
;
wire
CORETSE_AHBoI0I
;
wire
CORETSE_AHBiI0I
;
wire
CORETSE_AHBOl0I
;
wire
[
31
:
0
]
CORETSE_AHBIl0I
;
assign
CORETSE_AHBillI
=
CORETSE_AHBoi1
==
8
'h
12
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBiiOI
,
CORETSE_AHBOOII
,
CORETSE_AHBIOII
,
CORETSE_AHBlOII
,
CORETSE_AHBoOII
,
CORETSE_AHBioOI
,
CORETSE_AHBOiOI
,
CORETSE_AHBIiOI
,
CORETSE_AHBliOI
,
CORETSE_AHBoiOI
}
<=
#
CORETSE_AHBIoII
{
5
'h
00
,
5
'h
1F
}
;
else
if
(
CORETSE_AHBillI
)
{
CORETSE_AHBiiOI
,
CORETSE_AHBOOII
,
CORETSE_AHBIOII
,
CORETSE_AHBlOII
,
CORETSE_AHBoOII
,
CORETSE_AHBioOI
,
CORETSE_AHBOiOI
,
CORETSE_AHBIiOI
,
CORETSE_AHBliOI
,
CORETSE_AHBoiOI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
12
:
8
]
,
CORETSE_AHBii1
[
4
:
0
]
}
;
end
assign
CORETSE_AHBoolI
=
CORETSE_AHBoi1
==
8
'h
12
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBO0lI
=
CORETSE_AHBoi1
==
8
'h
13
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBi1OI
,
CORETSE_AHBl0OI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBIIlI
,
16
'h
FFFF
}
;
else
if
(
CORETSE_AHBO0lI
)
{
CORETSE_AHBi1OI
,
CORETSE_AHBl0OI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
(
RABITS
+
15
)
:
16
]
,
CORETSE_AHBii1
[
15
:
0
]
}
;
end
assign
CORETSE_AHBiolI
=
CORETSE_AHBoi1
==
8
'h
13
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBI0lI
=
CORETSE_AHBoi1
==
8
'h
14
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBo0OI
,
CORETSE_AHBi0OI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBIllI
,
CORETSE_AHBlllI
}
;
else
if
(
CORETSE_AHBI0lI
)
{
CORETSE_AHBo0OI
,
CORETSE_AHBi0OI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
(
RABITS
+
16
)
:
16
]
,
CORETSE_AHBii1
[
RABITS
:
0
]
}
;
end
assign
CORETSE_AHBOilI
=
CORETSE_AHBoi1
==
8
'h
14
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBl0lI
=
CORETSE_AHBoi1
==
8
'h
15
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBl1OI
,
CORETSE_AHBo1OI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBollI
,
CORETSE_AHBOIlI
}
;
else
if
(
CORETSE_AHBl0lI
)
{
CORETSE_AHBl1OI
,
CORETSE_AHBo1OI
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
(
TABITS
+
16
)
:
16
]
,
CORETSE_AHBii1
[
TABITS
:
0
]
}
;
end
assign
CORETSE_AHBIilI
=
CORETSE_AHBoi1
==
8
'h
15
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBo0lI
=
CORETSE_AHBoi1
==
8
'h
16
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBOoOI
[
17
:
0
]
<=
#
CORETSE_AHBIoII
18
'h
00008
;
else
if
(
CORETSE_AHBo0lI
)
CORETSE_AHBOoOI
[
17
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
17
:
0
]
;
end
assign
CORETSE_AHBlilI
=
CORETSE_AHBoi1
==
8
'h
16
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBi0lI
=
CORETSE_AHBoi1
==
8
'h
17
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBI1OI
,
CORETSE_AHBooOI
,
CORETSE_AHBO1OI
,
CORETSE_AHBloOI
,
CORETSE_AHBIoOI
[
17
:
0
]
}
<=
#
CORETSE_AHBIoII
22
'h
0B_FFF7
;
else
if
(
CORETSE_AHBi0lI
)
{
CORETSE_AHBI1OI
,
CORETSE_AHBooOI
,
CORETSE_AHBO1OI
,
CORETSE_AHBloOI
,
CORETSE_AHBIoOI
[
17
:
0
]
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
22
]
,
CORETSE_AHBii1
[
20
:
0
]
}
;
end
assign
CORETSE_AHBoilI
=
CORETSE_AHBoi1
==
8
'h
17
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBO1lI
=
CORETSE_AHBoi1
==
8
'h
18
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBOIII
,
CORETSE_AHBIIII
[
CORETSE_AHBIo1
+:
8
]
,
CORETSE_AHBiOII
}
<=
#
CORETSE_AHBIoII
{
9
'h
0
,
CORETSE_AHBlOlI
}
;
else
if
(
CORETSE_AHBO1lI
)
{
CORETSE_AHBOIII
,
CORETSE_AHBIIII
[
CORETSE_AHBIo1
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBiOII
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
]
,
CORETSE_AHBii1
[
16
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBii1
[
(
TABITS
+
1
)
:
0
]
}
;
end
assign
CORETSE_AHBiilI
=
CORETSE_AHBoi1
==
8
'h
18
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBI1lI
=
CORETSE_AHBoi1
==
8
'h
19
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBIIII
[
31
:
0
]
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
if
(
CORETSE_AHBI1lI
)
CORETSE_AHBIIII
[
31
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
31
:
0
]
;
end
assign
CORETSE_AHBOO0I
=
CORETSE_AHBoi1
==
8
'h
19
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
generate
if
(
CORETSE_AHBIo1
==
64
)
begin
assign
CORETSE_AHBl1lI
=
CORETSE_AHBoi1
==
8
'h
20
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBIIII
[
63
:
32
]
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
if
(
CORETSE_AHBl1lI
)
CORETSE_AHBIIII
[
63
:
32
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
31
:
0
]
;
end
assign
CORETSE_AHBIO0I
=
CORETSE_AHBoi1
==
8
'h
20
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
end
else
begin
assign
CORETSE_AHBIO0I
=
0
;
assign
CORETSE_AHBl1lI
=
0
;
end
endgenerate
assign
CORETSE_AHBo1lI
=
CORETSE_AHBoi1
==
8
'h
1a
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBoIII
,
CORETSE_AHBlIII
}
<=
#
CORETSE_AHBIoII
{
1
'b
0
,
CORETSE_AHBlOlI
}
;
else
if
(
CORETSE_AHBo1lI
)
{
CORETSE_AHBoIII
,
CORETSE_AHBlIII
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
]
,
CORETSE_AHBii1
[
(
TABITS
+
1
)
:
0
]
}
;
end
assign
CORETSE_AHBlO0I
=
CORETSE_AHBoi1
==
8
'h
1a
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBoO0I
=
CORETSE_AHBoi1
==
8
'h
1B
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
generate
if
(
CORETSE_AHBIo1
==
64
)
assign
CORETSE_AHBiO0I
=
CORETSE_AHBoi1
==
8
'h
21
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
else
assign
CORETSE_AHBiO0I
=
0
;
endgenerate
assign
CORETSE_AHBi1lI
=
CORETSE_AHBoi1
==
8
'h
1c
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBOlII
,
CORETSE_AHBIlII
[
CORETSE_AHBIo1
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBiIII
}
<=
#
CORETSE_AHBIoII
{
9
'h
0
,
CORETSE_AHBlIlI
}
;
else
if
(
CORETSE_AHBi1lI
)
{
CORETSE_AHBOlII
,
CORETSE_AHBIlII
[
CORETSE_AHBIo1
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBiIII
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
]
,
CORETSE_AHBii1
[
16
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBii1
[
RABITS
+
1
:
0
]
}
;
end
assign
CORETSE_AHBOI0I
=
CORETSE_AHBoi1
==
8
'h
1c
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBOolI
=
CORETSE_AHBoi1
==
8
'h
1d
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBIlII
[
31
:
0
]
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
if
(
CORETSE_AHBOolI
)
CORETSE_AHBIlII
[
31
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
31
:
0
]
;
end
assign
CORETSE_AHBII0I
=
CORETSE_AHBoi1
==
8
'h
1d
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
generate
if
(
CORETSE_AHBIo1
==
64
)
begin
assign
CORETSE_AHBIolI
=
CORETSE_AHBoi1
==
8
'h
22
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
CORETSE_AHBIlII
[
63
:
32
]
<=
#
CORETSE_AHBIoII
32
'h
0
;
else
if
(
CORETSE_AHBIolI
)
CORETSE_AHBIlII
[
63
:
32
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBii1
[
31
:
0
]
;
end
assign
CORETSE_AHBlI0I
=
CORETSE_AHBoi1
==
8
'h
22
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
end
else
begin
assign
CORETSE_AHBlI0I
=
0
;
assign
CORETSE_AHBll0I
=
0
;
end
endgenerate
assign
CORETSE_AHBlolI
=
CORETSE_AHBoi1
==
8
'h
1e
&
~
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
always
@
(
posedge
CORETSE_AHBOi1
or
posedge
CORETSE_AHBio1
)
begin
if
(
CORETSE_AHBio1
)
{
CORETSE_AHBolII
,
CORETSE_AHBllII
}
<=
#
CORETSE_AHBIoII
{
1
'b
0
,
CORETSE_AHBlIlI
}
;
else
if
(
CORETSE_AHBlolI
)
{
CORETSE_AHBolII
,
CORETSE_AHBllII
}
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBii1
[
31
]
,
CORETSE_AHBii1
[
RABITS
+
1
:
0
]
}
;
end
assign
CORETSE_AHBoI0I
=
CORETSE_AHBoi1
==
8
'h
1e
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBiI0I
=
CORETSE_AHBoi1
==
8
'h
1F
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
generate
if
(
CORETSE_AHBIo1
==
64
)
assign
CORETSE_AHBOl0I
=
CORETSE_AHBoi1
==
8
'h
23
&
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
else
assign
CORETSE_AHBOl0I
=
0
;
endgenerate
assign
CORETSE_AHBI1i
=
CORETSE_AHBli1
&
~
CORETSE_AHBIi1
;
assign
CORETSE_AHBO1i
=
{
32
{
CORETSE_AHBoolI
}
}
&
{
11
'h
0
,
CORETSE_AHBoOOI
,
CORETSE_AHBiOOI
,
CORETSE_AHBOIOI
,
CORETSE_AHBIIOI
,
CORETSE_AHBlIOI
,
3
'h
0
,
CORETSE_AHBiiOI
,
CORETSE_AHBOOII
,
CORETSE_AHBIOII
,
CORETSE_AHBlOII
,
CORETSE_AHBoOII
,
3
'h
0
,
CORETSE_AHBioOI
,
CORETSE_AHBOiOI
,
CORETSE_AHBIiOI
,
CORETSE_AHBliOI
,
CORETSE_AHBoiOI
}
|
{
32
{
CORETSE_AHBiolI
}
}
&
{
CORETSE_AHBoIlI
,
CORETSE_AHBi1OI
,
CORETSE_AHBl0OI
}
|
{
32
{
CORETSE_AHBOilI
}
}
&
{
CORETSE_AHBiIlI
,
CORETSE_AHBo0OI
,
CORETSE_AHBiIlI
,
CORETSE_AHBi0OI
}
|
{
32
{
CORETSE_AHBIilI
}
}
&
{
CORETSE_AHBoOlI
,
CORETSE_AHBl1OI
,
CORETSE_AHBoOlI
,
CORETSE_AHBo1OI
}
|
{
32
{
CORETSE_AHBlilI
}
}
&
{
14
'h
0
,
CORETSE_AHBOoOI
}
|
{
32
{
CORETSE_AHBoilI
}
}
&
{
9
'h
0
,
CORETSE_AHBI1OI
,
CORETSE_AHBoIOI
,
CORETSE_AHBooOI
,
CORETSE_AHBO1OI
,
CORETSE_AHBloOI
,
CORETSE_AHBIoOI
}
|
{
32
{
CORETSE_AHBiilI
}
}
&
{
CORETSE_AHBOIII
,
CORETSE_AHBiIOI
,
6
'h
0
,
CORETSE_AHBIIII
[
CORETSE_AHBIo1
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBoOlI
,
CORETSE_AHBOlOI
}
|
{
32
{
CORETSE_AHBOO0I
}
}
&
{
CORETSE_AHBIIII
[
31
:
0
]
}
|
{
32
{
CORETSE_AHBlO0I
}
}
&
{
CORETSE_AHBoIII
,
CORETSE_AHBIlOI
,
6
'h
0
,
CORETSE_AHBllOI
[
CORETSE_AHBIo1
+:
(
CORETSE_AHBlo1
+
6
)
]
,
16
'h
0000
}
|
{
32
{
CORETSE_AHBlO0I
}
}
&
{
CORETSE_AHBiOlI
,
CORETSE_AHBlIII
}
|
{
32
{
CORETSE_AHBoO0I
}
}
&
{
CORETSE_AHBllOI
[
31
:
0
]
}
|
{
32
{
CORETSE_AHBOI0I
}
}
&
{
CORETSE_AHBOlII
,
CORETSE_AHBolOI
,
6
'h
0
,
CORETSE_AHBIlII
[
(
CORETSE_AHBIo1
)
+:
(
CORETSE_AHBlo1
+
6
)
]
,
CORETSE_AHBiIlI
,
CORETSE_AHBilOI
}
|
{
32
{
CORETSE_AHBII0I
}
}
&
{
CORETSE_AHBIlII
[
31
:
0
]
}
|
{
32
{
CORETSE_AHBoI0I
}
}
&
{
CORETSE_AHBolII
,
CORETSE_AHBO0OI
,
6
'h
0
,
CORETSE_AHBI0OI
[
CORETSE_AHBIo1
+:
(
CORETSE_AHBlo1
+
6
)
]
,
{
{
16
-
RABITS
}
{
1
'h
0
}
}
,
CORETSE_AHBllII
}
|
{
32
{
CORETSE_AHBiI0I
}
}
&
{
CORETSE_AHBI0OI
[
31
:
0
]
}
|
CORETSE_AHBIl0I
;
generate
if
(
CORETSE_AHBIo1
==
64
)
begin
assign
CORETSE_AHBIl0I
=
{
32
{
CORETSE_AHBIO0I
}
}
&
{
CORETSE_AHBIIII
[
63
:
32
]
}
|
{
32
{
CORETSE_AHBiO0I
}
}
&
{
CORETSE_AHBllOI
[
63
:
32
]
}
|
{
32
{
CORETSE_AHBlI0I
}
}
&
{
CORETSE_AHBIlII
[
63
:
32
]
}
|
{
32
{
CORETSE_AHBOl0I
}
}
&
{
CORETSE_AHBI0OI
[
63
:
32
]
}
;
end
else
assign
CORETSE_AHBIl0I
=
32
'h
0
;
endgenerate
endmodule
