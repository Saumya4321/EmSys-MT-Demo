// REVISION    : $Revision: 1.2 $
//              Mentor Proprietary and Confidential
//              Copyright (c) 2000, Mentor Intellectual Property Development
`timescale 1ns/1ns
module
pemstat_eim
(
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
,
CORETSE_AHBliOi
,
CORETSE_AHBoiOi
,
CORETSE_AHBiiOi
,
CORETSE_AHBOOIi
,
CORETSE_AHBooOi
,
CORETSE_AHBioOi
,
CORETSE_AHBOlIi
,
CORETSE_AHBIlIi
,
CORETSE_AHBllIi
,
CORETSE_AHBolIi
,
CORETSE_AHBilIi
,
CORETSE_AHBO0Ii
,
CORETSE_AHBI0Ii
,
CORETSE_AHBl0Ii
,
CORETSE_AHBo0Ii
,
CORETSE_AHBi0Ii
,
CORETSE_AHBO1Ii
,
CORETSE_AHBI1Ii
,
CORETSE_AHBl1Ii
,
CORETSE_AHBo1Ii
,
CORETSE_AHBi1Ii
,
CORETSE_AHBOoIi
,
CORETSE_AHBIoIi
,
CORETSE_AHBloIi
,
CORETSE_AHBooIi
,
CORETSE_AHBioIi
,
CORETSE_AHBOiIi
,
CORETSE_AHBIiIi
,
CORETSE_AHBliIi
,
CORETSE_AHBoiIi
,
CORETSE_AHBiiIi
,
CORETSE_AHBOOli
,
CORETSE_AHBIOli
,
CORETSE_AHBlOli
,
CORETSE_AHBoOli
,
CORETSE_AHBiOli
,
CORETSE_AHBOIli
,
CORETSE_AHBIIli
,
CORETSE_AHBlIli
,
CORETSE_AHBoIli
,
CORETSE_AHBiIli
,
CORETSE_AHBOlli
,
CORETSE_AHBIlli
,
CORETSE_AHBllli
,
CORETSE_AHBolli
,
CORETSE_AHBilli
,
CORETSE_AHBO0li
,
CORETSE_AHBI0li
,
CORETSE_AHBl0li
,
CORETSE_AHBo0li
,
CORETSE_AHBi0li
,
CORETSE_AHBIOIi
,
CORETSE_AHBlOIi
,
CORETSE_AHBoOIi
,
CORETSE_AHBlIIi
,
CORETSE_AHBoIIi
,
CORETSE_AHBiIIi
)
;
input
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
;
input
[
6
:
0
]
CORETSE_AHBliOi
;
input
CORETSE_AHBoiOi
,
CORETSE_AHBiiOi
;
input
[
31
:
0
]
CORETSE_AHBOOIi
;
input
CORETSE_AHBooOi
,
CORETSE_AHBioOi
;
input
[
43
:
0
]
CORETSE_AHBOlIi
;
input
[
30
:
0
]
CORETSE_AHBIlIi
,
CORETSE_AHBllIi
,
CORETSE_AHBolIi
,
CORETSE_AHBilIi
,
CORETSE_AHBO0Ii
,
CORETSE_AHBI0Ii
,
CORETSE_AHBl0Ii
,
CORETSE_AHBo0Ii
;
input
[
30
:
0
]
CORETSE_AHBi0Ii
,
CORETSE_AHBO1Ii
,
CORETSE_AHBI1Ii
,
CORETSE_AHBl1Ii
,
CORETSE_AHBo1Ii
,
CORETSE_AHBi1Ii
,
CORETSE_AHBOoIi
,
CORETSE_AHBIoIi
;
input
[
30
:
0
]
CORETSE_AHBloIi
,
CORETSE_AHBooIi
,
CORETSE_AHBioIi
,
CORETSE_AHBOiIi
,
CORETSE_AHBIiIi
,
CORETSE_AHBliIi
,
CORETSE_AHBoiIi
,
CORETSE_AHBiiIi
;
input
[
30
:
0
]
CORETSE_AHBOOli
,
CORETSE_AHBIOli
,
CORETSE_AHBlOli
,
CORETSE_AHBoOli
,
CORETSE_AHBiOli
,
CORETSE_AHBOIli
,
CORETSE_AHBIIli
,
CORETSE_AHBlIli
;
input
[
30
:
0
]
CORETSE_AHBoIli
,
CORETSE_AHBiIli
,
CORETSE_AHBOlli
,
CORETSE_AHBIlli
,
CORETSE_AHBllli
,
CORETSE_AHBolli
,
CORETSE_AHBilli
,
CORETSE_AHBO0li
;
input
[
30
:
0
]
CORETSE_AHBI0li
,
CORETSE_AHBl0li
,
CORETSE_AHBo0li
,
CORETSE_AHBi0li
;
output
[
31
:
0
]
CORETSE_AHBIOIi
;
output
CORETSE_AHBlOIi
,
CORETSE_AHBoOIi
;
output
[
43
:
0
]
CORETSE_AHBlIIi
,
CORETSE_AHBoIIi
,
CORETSE_AHBiIIi
;
reg
CORETSE_AHBlOIi
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBlI0i
,
CORETSE_AHBoI0i
,
CORETSE_AHBiI0i
;
wire
CORETSE_AHBOl0i
;
reg
CORETSE_AHBIl0i
,
CORETSE_AHBll0i
,
CORETSE_AHBol0i
;
wire
CORETSE_AHBil0i
;
wire
[
43
:
0
]
CORETSE_AHBO00i
;
wire
[
30
:
0
]
CORETSE_AHBI00i
;
reg
[
30
:
0
]
CORETSE_AHBl00i
;
wire
CORETSE_AHBo00i
,
CORETSE_AHBi00i
,
CORETSE_AHBO10i
,
CORETSE_AHBI10i
;
reg
[
23
:
0
]
CORETSE_AHBl10i
;
reg
[
19
:
0
]
CORETSE_AHBo10i
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBlI0i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlI0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiOi
;
end
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBoI0i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoI0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBlI0i
;
end
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBiI0i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiI0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI0i
;
end
assign
CORETSE_AHBOl0i
=
CORETSE_AHBoI0i
&
~
CORETSE_AHBiI0i
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBlOIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBlOIi
&
~
CORETSE_AHBoI0i
)
CORETSE_AHBlOIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
~
CORETSE_AHBlOIi
&
CORETSE_AHBoI0i
&
~
CORETSE_AHBiiOi
&
(
CORETSE_AHBliOi
>=
7
'h
20
)
&
(
CORETSE_AHBliOi
<=
7
'h
5F
)
)
CORETSE_AHBlOIi
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
~
CORETSE_AHBlOIi
&
CORETSE_AHBiI0i
&
CORETSE_AHBiiOi
&
(
CORETSE_AHBliOi
>=
7
'h
20
)
&
(
CORETSE_AHBliOi
<=
7
'h
5F
)
)
CORETSE_AHBlOIi
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBIl0i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIl0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBioOi
;
end
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBll0i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBll0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl0i
;
end
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBol0i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBol0i
<=
#
CORETSE_AHBIoII
CORETSE_AHBll0i
;
end
assign
CORETSE_AHBil0i
=
CORETSE_AHBll0i
&
~
CORETSE_AHBol0i
;
assign
CORETSE_AHBO00i
[
00
]
=
(
CORETSE_AHBliOi
==
7
'h
20
)
;
assign
CORETSE_AHBO00i
[
01
]
=
(
CORETSE_AHBliOi
==
7
'h
21
)
;
assign
CORETSE_AHBO00i
[
02
]
=
(
CORETSE_AHBliOi
==
7
'h
22
)
;
assign
CORETSE_AHBO00i
[
03
]
=
(
CORETSE_AHBliOi
==
7
'h
23
)
;
assign
CORETSE_AHBO00i
[
04
]
=
(
CORETSE_AHBliOi
==
7
'h
24
)
;
assign
CORETSE_AHBO00i
[
05
]
=
(
CORETSE_AHBliOi
==
7
'h
25
)
;
assign
CORETSE_AHBO00i
[
06
]
=
(
CORETSE_AHBliOi
==
7
'h
26
)
;
assign
CORETSE_AHBO00i
[
07
]
=
(
CORETSE_AHBliOi
==
7
'h
27
)
;
assign
CORETSE_AHBO00i
[
08
]
=
(
CORETSE_AHBliOi
==
7
'h
28
)
;
assign
CORETSE_AHBO00i
[
09
]
=
(
CORETSE_AHBliOi
==
7
'h
29
)
;
assign
CORETSE_AHBO00i
[
10
]
=
(
CORETSE_AHBliOi
==
7
'h
2A
)
;
assign
CORETSE_AHBO00i
[
11
]
=
(
CORETSE_AHBliOi
==
7
'h
2B
)
;
assign
CORETSE_AHBO00i
[
12
]
=
(
CORETSE_AHBliOi
==
7
'h
2C
)
;
assign
CORETSE_AHBO00i
[
13
]
=
(
CORETSE_AHBliOi
==
7
'h
2D
)
;
assign
CORETSE_AHBO00i
[
14
]
=
(
CORETSE_AHBliOi
==
7
'h
2E
)
;
assign
CORETSE_AHBO00i
[
15
]
=
(
CORETSE_AHBliOi
==
7
'h
2F
)
;
assign
CORETSE_AHBO00i
[
16
]
=
(
CORETSE_AHBliOi
==
7
'h
30
)
;
assign
CORETSE_AHBO00i
[
17
]
=
(
CORETSE_AHBliOi
==
7
'h
31
)
;
assign
CORETSE_AHBO00i
[
18
]
=
(
CORETSE_AHBliOi
==
7
'h
32
)
;
assign
CORETSE_AHBO00i
[
19
]
=
(
CORETSE_AHBliOi
==
7
'h
33
)
;
assign
CORETSE_AHBO00i
[
20
]
=
(
CORETSE_AHBliOi
==
7
'h
34
)
;
assign
CORETSE_AHBO00i
[
21
]
=
(
CORETSE_AHBliOi
==
7
'h
35
)
;
assign
CORETSE_AHBO00i
[
22
]
=
(
CORETSE_AHBliOi
==
7
'h
36
)
;
assign
CORETSE_AHBO00i
[
23
]
=
(
CORETSE_AHBliOi
==
7
'h
37
)
;
assign
CORETSE_AHBO00i
[
24
]
=
(
CORETSE_AHBliOi
==
7
'h
38
)
;
assign
CORETSE_AHBO00i
[
25
]
=
(
CORETSE_AHBliOi
==
7
'h
39
)
;
assign
CORETSE_AHBO00i
[
26
]
=
(
CORETSE_AHBliOi
==
7
'h
3A
)
;
assign
CORETSE_AHBO00i
[
27
]
=
(
CORETSE_AHBliOi
==
7
'h
3B
)
;
assign
CORETSE_AHBO00i
[
28
]
=
(
CORETSE_AHBliOi
==
7
'h
3C
)
;
assign
CORETSE_AHBO00i
[
29
]
=
(
CORETSE_AHBliOi
==
7
'h
3D
)
;
assign
CORETSE_AHBO00i
[
30
]
=
(
CORETSE_AHBliOi
==
7
'h
3E
)
;
assign
CORETSE_AHBO00i
[
31
]
=
(
CORETSE_AHBliOi
==
7
'h
3F
)
;
assign
CORETSE_AHBO00i
[
32
]
=
(
CORETSE_AHBliOi
==
7
'h
40
)
;
assign
CORETSE_AHBO00i
[
33
]
=
(
CORETSE_AHBliOi
==
7
'h
41
)
;
assign
CORETSE_AHBO00i
[
34
]
=
(
CORETSE_AHBliOi
==
7
'h
42
)
;
assign
CORETSE_AHBO00i
[
35
]
=
(
CORETSE_AHBliOi
==
7
'h
43
)
;
assign
CORETSE_AHBO00i
[
36
]
=
(
CORETSE_AHBliOi
==
7
'h
44
)
;
assign
CORETSE_AHBO00i
[
37
]
=
(
CORETSE_AHBliOi
==
7
'h
45
)
;
assign
CORETSE_AHBO00i
[
38
]
=
(
CORETSE_AHBliOi
==
7
'h
46
)
;
assign
CORETSE_AHBO00i
[
39
]
=
(
CORETSE_AHBliOi
==
7
'h
47
)
;
assign
CORETSE_AHBO00i
[
40
]
=
(
CORETSE_AHBliOi
==
7
'h
48
)
;
assign
CORETSE_AHBO00i
[
41
]
=
(
CORETSE_AHBliOi
==
7
'h
49
)
;
assign
CORETSE_AHBO00i
[
42
]
=
(
CORETSE_AHBliOi
==
7
'h
4A
)
;
assign
CORETSE_AHBO00i
[
43
]
=
(
CORETSE_AHBliOi
==
7
'h
4B
)
;
assign
CORETSE_AHBI00i
=
{
31
{
CORETSE_AHBO00i
[
00
]
}
}
&
{
CORETSE_AHBIlIi
}
|
{
31
{
CORETSE_AHBO00i
[
01
]
}
}
&
{
CORETSE_AHBllIi
}
|
{
31
{
CORETSE_AHBO00i
[
02
]
}
}
&
{
CORETSE_AHBolIi
}
|
{
31
{
CORETSE_AHBO00i
[
03
]
}
}
&
{
CORETSE_AHBilIi
}
|
{
31
{
CORETSE_AHBO00i
[
04
]
}
}
&
{
CORETSE_AHBO0Ii
}
|
{
31
{
CORETSE_AHBO00i
[
05
]
}
}
&
{
CORETSE_AHBI0Ii
}
|
{
31
{
CORETSE_AHBO00i
[
06
]
}
}
&
{
CORETSE_AHBl0Ii
}
|
{
31
{
CORETSE_AHBO00i
[
07
]
}
}
&
{
CORETSE_AHBo0Ii
}
|
{
31
{
CORETSE_AHBO00i
[
08
]
}
}
&
{
CORETSE_AHBi0Ii
}
|
{
31
{
CORETSE_AHBO00i
[
09
]
}
}
&
{
CORETSE_AHBO1Ii
}
|
{
31
{
CORETSE_AHBO00i
[
10
]
}
}
&
{
CORETSE_AHBI1Ii
}
|
{
31
{
CORETSE_AHBO00i
[
11
]
}
}
&
{
CORETSE_AHBl1Ii
}
|
{
31
{
CORETSE_AHBO00i
[
12
]
}
}
&
{
CORETSE_AHBo1Ii
}
|
{
31
{
CORETSE_AHBO00i
[
13
]
}
}
&
{
CORETSE_AHBi1Ii
}
|
{
31
{
CORETSE_AHBO00i
[
14
]
}
}
&
{
CORETSE_AHBOoIi
}
|
{
31
{
CORETSE_AHBO00i
[
15
]
}
}
&
{
CORETSE_AHBIoIi
}
|
{
31
{
CORETSE_AHBO00i
[
16
]
}
}
&
{
CORETSE_AHBloIi
}
|
{
31
{
CORETSE_AHBO00i
[
17
]
}
}
&
{
CORETSE_AHBooIi
}
|
{
31
{
CORETSE_AHBO00i
[
18
]
}
}
&
{
CORETSE_AHBioIi
}
|
{
31
{
CORETSE_AHBO00i
[
19
]
}
}
&
{
CORETSE_AHBOiIi
}
|
{
31
{
CORETSE_AHBO00i
[
20
]
}
}
&
{
CORETSE_AHBIiIi
}
|
{
31
{
CORETSE_AHBO00i
[
21
]
}
}
&
{
CORETSE_AHBliIi
}
|
{
31
{
CORETSE_AHBO00i
[
22
]
}
}
&
{
CORETSE_AHBoiIi
}
|
{
31
{
CORETSE_AHBO00i
[
23
]
}
}
&
{
CORETSE_AHBiiIi
}
|
{
31
{
CORETSE_AHBO00i
[
24
]
}
}
&
{
CORETSE_AHBOOli
}
|
{
31
{
CORETSE_AHBO00i
[
25
]
}
}
&
{
CORETSE_AHBIOli
}
|
{
31
{
CORETSE_AHBO00i
[
26
]
}
}
&
{
CORETSE_AHBlOli
}
|
{
31
{
CORETSE_AHBO00i
[
27
]
}
}
&
{
CORETSE_AHBoOli
}
|
{
31
{
CORETSE_AHBO00i
[
28
]
}
}
&
{
CORETSE_AHBiOli
}
|
{
31
{
CORETSE_AHBO00i
[
29
]
}
}
&
{
CORETSE_AHBOIli
}
|
{
31
{
CORETSE_AHBO00i
[
30
]
}
}
&
{
CORETSE_AHBIIli
}
|
{
31
{
CORETSE_AHBO00i
[
31
]
}
}
&
{
CORETSE_AHBlIli
}
|
{
31
{
CORETSE_AHBO00i
[
32
]
}
}
&
{
CORETSE_AHBoIli
}
|
{
31
{
CORETSE_AHBO00i
[
33
]
}
}
&
{
CORETSE_AHBiIli
}
|
{
31
{
CORETSE_AHBO00i
[
34
]
}
}
&
{
CORETSE_AHBOlli
}
|
{
31
{
CORETSE_AHBO00i
[
35
]
}
}
&
{
CORETSE_AHBIlli
}
|
{
31
{
CORETSE_AHBO00i
[
36
]
}
}
&
{
CORETSE_AHBllli
}
|
{
31
{
CORETSE_AHBO00i
[
37
]
}
}
&
{
CORETSE_AHBolli
}
|
{
31
{
CORETSE_AHBO00i
[
38
]
}
}
&
{
CORETSE_AHBilli
}
|
{
31
{
CORETSE_AHBO00i
[
39
]
}
}
&
{
CORETSE_AHBO0li
}
|
{
31
{
CORETSE_AHBO00i
[
40
]
}
}
&
{
CORETSE_AHBI0li
}
|
{
31
{
CORETSE_AHBO00i
[
41
]
}
}
&
{
CORETSE_AHBl0li
}
|
{
31
{
CORETSE_AHBO00i
[
42
]
}
}
&
{
CORETSE_AHBo0li
}
|
{
31
{
CORETSE_AHBO00i
[
43
]
}
}
&
{
CORETSE_AHBi0li
}
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBl00i
<=
#
CORETSE_AHBIoII
31
'h
0
;
else
if
(
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
CORETSE_AHBl00i
<=
#
CORETSE_AHBIoII
CORETSE_AHBI00i
;
end
assign
CORETSE_AHBo00i
=
(
CORETSE_AHBliOi
==
7
'h
4C
)
&
CORETSE_AHBoI0i
;
assign
CORETSE_AHBi00i
=
(
CORETSE_AHBliOi
==
7
'h
4D
)
&
CORETSE_AHBoI0i
;
assign
CORETSE_AHBO10i
=
(
CORETSE_AHBliOi
==
7
'h
4E
)
&
CORETSE_AHBoI0i
;
assign
CORETSE_AHBI10i
=
(
CORETSE_AHBliOi
==
7
'h
4F
)
&
CORETSE_AHBoI0i
;
assign
CORETSE_AHBIOIi
=
{
32
{
(
|
CORETSE_AHBO00i
&
CORETSE_AHBoI0i
&
CORETSE_AHBiiOi
)
}
}
&
{
1
'b
0
,
CORETSE_AHBl00i
}
|
{
32
{
(
CORETSE_AHBo00i
&
CORETSE_AHBoI0i
&
CORETSE_AHBiiOi
)
}
}
&
{
CORETSE_AHBOlIi
[
0
]
,
CORETSE_AHBOlIi
[
1
]
,
CORETSE_AHBOlIi
[
2
]
,
CORETSE_AHBOlIi
[
3
]
,
CORETSE_AHBOlIi
[
4
]
,
CORETSE_AHBOlIi
[
5
]
,
CORETSE_AHBOlIi
[
6
]
,
1
'h
0
,
4
'h
0
,
3
'h
0
,
CORETSE_AHBOlIi
[
7
]
,
CORETSE_AHBOlIi
[
8
]
,
CORETSE_AHBOlIi
[
9
]
,
CORETSE_AHBOlIi
[
10
]
,
CORETSE_AHBOlIi
[
11
]
,
CORETSE_AHBOlIi
[
12
]
,
CORETSE_AHBOlIi
[
13
]
,
CORETSE_AHBOlIi
[
14
]
,
CORETSE_AHBOlIi
[
15
]
,
CORETSE_AHBOlIi
[
16
]
,
CORETSE_AHBOlIi
[
17
]
,
CORETSE_AHBOlIi
[
18
]
,
CORETSE_AHBOlIi
[
19
]
,
CORETSE_AHBOlIi
[
20
]
,
CORETSE_AHBOlIi
[
21
]
,
CORETSE_AHBOlIi
[
22
]
,
CORETSE_AHBOlIi
[
23
]
}
|
{
32
{
(
CORETSE_AHBi00i
&
CORETSE_AHBoI0i
&
CORETSE_AHBiiOi
)
}
}
&
{
12
'h
0
,
CORETSE_AHBOlIi
[
38
]
,
CORETSE_AHBOlIi
[
39
]
,
CORETSE_AHBOlIi
[
40
]
,
CORETSE_AHBOlIi
[
41
]
,
CORETSE_AHBOlIi
[
42
]
,
CORETSE_AHBOlIi
[
43
]
,
CORETSE_AHBOlIi
[
24
]
,
CORETSE_AHBOlIi
[
25
]
,
CORETSE_AHBOlIi
[
26
]
,
CORETSE_AHBOlIi
[
27
]
,
CORETSE_AHBOlIi
[
28
]
,
CORETSE_AHBOlIi
[
29
]
,
CORETSE_AHBOlIi
[
30
]
,
CORETSE_AHBOlIi
[
31
]
,
CORETSE_AHBOlIi
[
32
]
,
CORETSE_AHBOlIi
[
33
]
,
CORETSE_AHBOlIi
[
34
]
,
CORETSE_AHBOlIi
[
35
]
,
CORETSE_AHBOlIi
[
36
]
,
CORETSE_AHBOlIi
[
37
]
}
|
{
32
{
(
CORETSE_AHBO10i
&
CORETSE_AHBoI0i
&
CORETSE_AHBiiOi
)
}
}
&
{
CORETSE_AHBl10i
[
23
:
17
]
,
8
'h
0
,
CORETSE_AHBl10i
[
16
:
0
]
}
|
{
32
{
(
CORETSE_AHBI10i
&
CORETSE_AHBoI0i
&
CORETSE_AHBiiOi
)
}
}
&
{
12
'h
0
,
CORETSE_AHBo10i
[
19
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBl10i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
24
'h
FFFFFF
;
else
if
(
CORETSE_AHBO10i
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
CORETSE_AHBl10i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBOOIi
[
31
:
25
]
,
CORETSE_AHBOOIi
[
16
:
0
]
}
;
end
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBo10i
[
19
:
0
]
<=
#
CORETSE_AHBIoII
20
'h
FFFFF
;
else
if
(
CORETSE_AHBI10i
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
CORETSE_AHBo10i
[
19
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOIi
[
19
:
0
]
;
end
assign
CORETSE_AHBoOIi
=
|
(
CORETSE_AHBOlIi
&
~
{
CORETSE_AHBo10i
[
14
]
,
CORETSE_AHBo10i
[
15
]
,
CORETSE_AHBo10i
[
16
]
,
CORETSE_AHBo10i
[
17
]
,
CORETSE_AHBo10i
[
18
]
,
CORETSE_AHBo10i
[
19
]
,
CORETSE_AHBo10i
[
0
]
,
CORETSE_AHBo10i
[
1
]
,
CORETSE_AHBo10i
[
2
]
,
CORETSE_AHBo10i
[
3
]
,
CORETSE_AHBo10i
[
4
]
,
CORETSE_AHBo10i
[
5
]
,
CORETSE_AHBo10i
[
6
]
,
CORETSE_AHBo10i
[
7
]
,
CORETSE_AHBo10i
[
8
]
,
CORETSE_AHBo10i
[
9
]
,
CORETSE_AHBo10i
[
10
]
,
CORETSE_AHBo10i
[
11
]
,
CORETSE_AHBo10i
[
12
]
,
CORETSE_AHBo10i
[
13
]
,
CORETSE_AHBl10i
[
0
]
,
CORETSE_AHBl10i
[
1
]
,
CORETSE_AHBl10i
[
2
]
,
CORETSE_AHBl10i
[
3
]
,
CORETSE_AHBl10i
[
4
]
,
CORETSE_AHBl10i
[
5
]
,
CORETSE_AHBl10i
[
6
]
,
CORETSE_AHBl10i
[
7
]
,
CORETSE_AHBl10i
[
8
]
,
CORETSE_AHBl10i
[
9
]
,
CORETSE_AHBl10i
[
10
]
,
CORETSE_AHBl10i
[
11
]
,
CORETSE_AHBl10i
[
12
]
,
CORETSE_AHBl10i
[
13
]
,
CORETSE_AHBl10i
[
14
]
,
CORETSE_AHBl10i
[
15
]
,
CORETSE_AHBl10i
[
16
]
,
CORETSE_AHBl10i
[
17
]
,
CORETSE_AHBl10i
[
18
]
,
CORETSE_AHBl10i
[
19
]
,
CORETSE_AHBl10i
[
20
]
,
CORETSE_AHBl10i
[
21
]
,
CORETSE_AHBl10i
[
22
]
,
CORETSE_AHBl10i
[
23
]
}
)
;
assign
CORETSE_AHBiIIi
[
23
:
0
]
=
{
24
{
(
CORETSE_AHBo00i
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
}
}
&
{
CORETSE_AHBOOIi
[
0
]
,
CORETSE_AHBOOIi
[
1
]
,
CORETSE_AHBOOIi
[
2
]
,
CORETSE_AHBOOIi
[
3
]
,
CORETSE_AHBOOIi
[
4
]
,
CORETSE_AHBOOIi
[
5
]
,
CORETSE_AHBOOIi
[
6
]
,
CORETSE_AHBOOIi
[
7
]
,
CORETSE_AHBOOIi
[
8
]
,
CORETSE_AHBOOIi
[
9
]
,
CORETSE_AHBOOIi
[
10
]
,
CORETSE_AHBOOIi
[
11
]
,
CORETSE_AHBOOIi
[
12
]
,
CORETSE_AHBOOIi
[
13
]
,
CORETSE_AHBOOIi
[
14
]
,
CORETSE_AHBOOIi
[
15
]
,
CORETSE_AHBOOIi
[
16
]
,
CORETSE_AHBOOIi
[
25
]
,
CORETSE_AHBOOIi
[
26
]
,
CORETSE_AHBOOIi
[
27
]
,
CORETSE_AHBOOIi
[
28
]
,
CORETSE_AHBOOIi
[
29
]
,
CORETSE_AHBOOIi
[
30
]
,
CORETSE_AHBOOIi
[
31
]
}
;
assign
CORETSE_AHBiIIi
[
43
:
24
]
=
{
20
{
(
CORETSE_AHBi00i
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
}
}
&
{
CORETSE_AHBOOIi
[
14
]
,
CORETSE_AHBOOIi
[
15
]
,
CORETSE_AHBOOIi
[
16
]
,
CORETSE_AHBOOIi
[
17
]
,
CORETSE_AHBOOIi
[
18
]
,
CORETSE_AHBOOIi
[
19
]
,
CORETSE_AHBOOIi
[
0
]
,
CORETSE_AHBOOIi
[
1
]
,
CORETSE_AHBOOIi
[
2
]
,
CORETSE_AHBOOIi
[
3
]
,
CORETSE_AHBOOIi
[
4
]
,
CORETSE_AHBOOIi
[
5
]
,
CORETSE_AHBOOIi
[
6
]
,
CORETSE_AHBOOIi
[
7
]
,
CORETSE_AHBOOIi
[
8
]
,
CORETSE_AHBOOIi
[
9
]
,
CORETSE_AHBOOIi
[
10
]
,
CORETSE_AHBOOIi
[
11
]
,
CORETSE_AHBOOIi
[
12
]
,
CORETSE_AHBOOIi
[
13
]
}
;
assign
CORETSE_AHBlIIi
[
00
]
=
(
CORETSE_AHBO00i
[
00
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
01
]
=
(
CORETSE_AHBO00i
[
01
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
02
]
=
(
CORETSE_AHBO00i
[
02
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
03
]
=
(
CORETSE_AHBO00i
[
03
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
04
]
=
(
CORETSE_AHBO00i
[
04
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
05
]
=
(
CORETSE_AHBO00i
[
05
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
06
]
=
(
CORETSE_AHBO00i
[
06
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
07
]
=
(
CORETSE_AHBO00i
[
07
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
08
]
=
(
CORETSE_AHBO00i
[
08
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
09
]
=
(
CORETSE_AHBO00i
[
09
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
10
]
=
(
CORETSE_AHBO00i
[
10
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
11
]
=
(
CORETSE_AHBO00i
[
11
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
12
]
=
(
CORETSE_AHBO00i
[
12
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
13
]
=
(
CORETSE_AHBO00i
[
13
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
14
]
=
(
CORETSE_AHBO00i
[
14
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
15
]
=
(
CORETSE_AHBO00i
[
15
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
16
]
=
(
CORETSE_AHBO00i
[
16
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
17
]
=
(
CORETSE_AHBO00i
[
17
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
18
]
=
(
CORETSE_AHBO00i
[
18
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
19
]
=
(
CORETSE_AHBO00i
[
19
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
20
]
=
(
CORETSE_AHBO00i
[
20
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
21
]
=
(
CORETSE_AHBO00i
[
21
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
22
]
=
(
CORETSE_AHBO00i
[
22
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
23
]
=
(
CORETSE_AHBO00i
[
23
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
24
]
=
(
CORETSE_AHBO00i
[
24
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
25
]
=
(
CORETSE_AHBO00i
[
25
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
26
]
=
(
CORETSE_AHBO00i
[
26
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
27
]
=
(
CORETSE_AHBO00i
[
27
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
28
]
=
(
CORETSE_AHBO00i
[
28
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
29
]
=
(
CORETSE_AHBO00i
[
29
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
30
]
=
(
CORETSE_AHBO00i
[
30
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
31
]
=
(
CORETSE_AHBO00i
[
31
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
32
]
=
(
CORETSE_AHBO00i
[
32
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
33
]
=
(
CORETSE_AHBO00i
[
33
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
34
]
=
(
CORETSE_AHBO00i
[
34
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
35
]
=
(
CORETSE_AHBO00i
[
35
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
36
]
=
(
CORETSE_AHBO00i
[
36
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
37
]
=
(
CORETSE_AHBO00i
[
37
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
38
]
=
(
CORETSE_AHBO00i
[
38
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
39
]
=
(
CORETSE_AHBO00i
[
39
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
40
]
=
(
CORETSE_AHBO00i
[
40
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
41
]
=
(
CORETSE_AHBO00i
[
41
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
42
]
=
(
CORETSE_AHBO00i
[
42
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBlIIi
[
43
]
=
(
CORETSE_AHBO00i
[
43
]
&
CORETSE_AHBooOi
&
CORETSE_AHBOl0i
&
CORETSE_AHBiiOi
)
|
CORETSE_AHBil0i
;
assign
CORETSE_AHBoIIi
[
00
]
=
(
CORETSE_AHBO00i
[
00
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
01
]
=
(
CORETSE_AHBO00i
[
01
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
02
]
=
(
CORETSE_AHBO00i
[
02
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
03
]
=
(
CORETSE_AHBO00i
[
03
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
04
]
=
(
CORETSE_AHBO00i
[
04
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
05
]
=
(
CORETSE_AHBO00i
[
05
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
06
]
=
(
CORETSE_AHBO00i
[
06
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
07
]
=
(
CORETSE_AHBO00i
[
07
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
08
]
=
(
CORETSE_AHBO00i
[
08
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
09
]
=
(
CORETSE_AHBO00i
[
09
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
10
]
=
(
CORETSE_AHBO00i
[
10
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
11
]
=
(
CORETSE_AHBO00i
[
11
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
12
]
=
(
CORETSE_AHBO00i
[
12
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
13
]
=
(
CORETSE_AHBO00i
[
13
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
14
]
=
(
CORETSE_AHBO00i
[
14
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
15
]
=
(
CORETSE_AHBO00i
[
15
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
16
]
=
(
CORETSE_AHBO00i
[
16
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
17
]
=
(
CORETSE_AHBO00i
[
17
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
18
]
=
(
CORETSE_AHBO00i
[
18
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
19
]
=
(
CORETSE_AHBO00i
[
19
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
20
]
=
(
CORETSE_AHBO00i
[
20
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
21
]
=
(
CORETSE_AHBO00i
[
21
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
22
]
=
(
CORETSE_AHBO00i
[
22
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
23
]
=
(
CORETSE_AHBO00i
[
23
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
24
]
=
(
CORETSE_AHBO00i
[
24
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
25
]
=
(
CORETSE_AHBO00i
[
25
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
26
]
=
(
CORETSE_AHBO00i
[
26
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
27
]
=
(
CORETSE_AHBO00i
[
27
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
28
]
=
(
CORETSE_AHBO00i
[
28
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
29
]
=
(
CORETSE_AHBO00i
[
29
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
30
]
=
(
CORETSE_AHBO00i
[
30
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
31
]
=
(
CORETSE_AHBO00i
[
31
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
32
]
=
(
CORETSE_AHBO00i
[
32
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
33
]
=
(
CORETSE_AHBO00i
[
33
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
34
]
=
(
CORETSE_AHBO00i
[
34
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
35
]
=
(
CORETSE_AHBO00i
[
35
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
36
]
=
(
CORETSE_AHBO00i
[
36
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
37
]
=
(
CORETSE_AHBO00i
[
37
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
38
]
=
(
CORETSE_AHBO00i
[
38
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
39
]
=
(
CORETSE_AHBO00i
[
39
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
40
]
=
(
CORETSE_AHBO00i
[
40
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
41
]
=
(
CORETSE_AHBO00i
[
41
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
42
]
=
(
CORETSE_AHBO00i
[
42
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
assign
CORETSE_AHBoIIi
[
43
]
=
(
CORETSE_AHBO00i
[
43
]
&
CORETSE_AHBOl0i
&
~
CORETSE_AHBiiOi
)
;
endmodule
