// REVISION    : $Revision: 1.12 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxrfif_sys
#
(
parameter
CORETSE_AHBoOI
=
0
,
parameter
RABITS
=
12
,
parameter
CORETSE_AHBIo1
=
32
,
parameter
CORETSE_AHBlo1
=
$clog2
(
CORETSE_AHBIo1
/
8
)
)
(
CORETSE_AHBii0
,
CORETSE_AHBl0o
,
CORETSE_AHBl0II
,
CORETSE_AHBlOII
,
CORETSE_AHBi1OI
,
CORETSE_AHBOoOI
,
CORETSE_AHBIoOI
,
CORETSE_AHBloOI
,
CORETSE_AHBooOI
,
CORETSE_AHBo0o
,
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
,
CORETSE_AHBl1o
,
CORETSE_AHBo1o
,
CORETSE_AHBi1o
,
CORETSE_AHBOoo
,
CORETSE_AHBooi
,
CORETSE_AHBlOOI
,
CORETSE_AHBioi
,
CORETSE_AHBOii
,
CORETSE_AHBiIII
,
CORETSE_AHBOlII
,
CORETSE_AHBIlII
,
CORETSE_AHBIIOI
,
CORETSE_AHBoIOI
,
CORETSE_AHBI0i
,
CORETSE_AHBl0i
,
CORETSE_AHBO0i
,
CORETSE_AHBIii
,
CORETSE_AHBlii
,
CORETSE_AHBiii
,
CORETSE_AHBOOOI
,
CORETSE_AHBIOOI
,
CORETSE_AHBoii
,
CORETSE_AHBolOI
,
CORETSE_AHBilOI
)
;
input
CORETSE_AHBii0
;
input
CORETSE_AHBl0o
;
input
CORETSE_AHBl0II
;
input
CORETSE_AHBlOII
;
input
[
RABITS
-
1
:
0
]
CORETSE_AHBi1OI
;
input
[
17
:
0
]
CORETSE_AHBOoOI
;
input
[
17
:
0
]
CORETSE_AHBIoOI
;
input
CORETSE_AHBloOI
;
input
CORETSE_AHBooOI
;
input
[
7
:
0
]
CORETSE_AHBo0o
;
input
CORETSE_AHBi0o
;
input
CORETSE_AHBO1o
;
input
CORETSE_AHBI1o
;
input
[
32
:
0
]
CORETSE_AHBl1o
;
input
CORETSE_AHBo1o
;
input
CORETSE_AHBi1o
;
input
CORETSE_AHBOoo
;
input
CORETSE_AHBooi
;
input
CORETSE_AHBlOOI
;
input
[
RABITS
:
0
]
CORETSE_AHBioi
;
input
CORETSE_AHBOii
;
input
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBiIII
;
input
CORETSE_AHBOlII
;
input
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIlII
;
output
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBI0i
;
output
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBl0i
;
output
CORETSE_AHBO0i
;
output
CORETSE_AHBIIOI
;
output
CORETSE_AHBoIOI
;
output
[
RABITS
:
0
]
CORETSE_AHBIii
;
output
CORETSE_AHBlii
;
output
[
RABITS
:
0
]
CORETSE_AHBiii
;
output
[
RABITS
:
0
]
CORETSE_AHBOOOI
;
output
CORETSE_AHBIOOI
;
output
CORETSE_AHBoii
;
output
CORETSE_AHBolOI
;
output
[
RABITS
:
0
]
CORETSE_AHBilOI
;
parameter
CORETSE_AHBlO1I
=
{
(
RABITS
+
2
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBoO1I
=
{
(
RABITS
+
1
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBol0I
=
{
(
RABITS
+
CORETSE_AHBlo1
+
1
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBIoII
=
1
;
wire
[
(
RABITS
+
CORETSE_AHBlo1
)
:
0
]
CORETSE_AHBiO1I
;
reg
[
(
RABITS
+
CORETSE_AHBlo1
)
:
0
]
CORETSE_AHBOI1I
,
CORETSE_AHBII1I
;
reg
CORETSE_AHBlI1I
;
wire
CORETSE_AHBoI1I
;
reg
CORETSE_AHBiI1I
,
CORETSE_AHBOl1I
;
wire
[
(
RABITS
+
CORETSE_AHBlo1
)
:
0
]
CORETSE_AHBIl1I
,
CORETSE_AHBll1I
;
reg
CORETSE_AHBol1I
;
reg
CORETSE_AHBIIOI
;
reg
[
RABITS
:
0
]
CORETSE_AHBIii
,
CORETSE_AHBiii
,
CORETSE_AHBOOOI
,
CORETSE_AHBil1I
;
reg
CORETSE_AHBlii
,
CORETSE_AHBIOOI
;
reg
CORETSE_AHBoii
;
wire
CORETSE_AHBO01I
;
reg
CORETSE_AHBI01I
;
reg
CORETSE_AHBoIOI
;
reg
CORETSE_AHBl01I
,
CORETSE_AHBo01I
;
reg
[
RABITS
:
0
]
CORETSE_AHBi01I
;
reg
CORETSE_AHBO11I
,
CORETSE_AHBI11I
;
reg
CORETSE_AHBl11I
,
CORETSE_AHBo11I
;
reg
CORETSE_AHBi11I
,
CORETSE_AHBOo1I
;
reg
CORETSE_AHBIo1I
,
CORETSE_AHBlo1I
;
wire
CORETSE_AHBoo1I
,
CORETSE_AHBio1I
;
reg
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBl0i
;
reg
CORETSE_AHBOi1I
;
reg
[
(
RABITS
+
CORETSE_AHBlo1
)
-
1
:
0
]
CORETSE_AHBIi1I
;
reg
CORETSE_AHBli1I
;
reg
CORETSE_AHBoi1I
;
reg
CORETSE_AHBii1I
;
wire
CORETSE_AHBOOoI
;
wire
CORETSE_AHBIOoI
;
wire
CORETSE_AHBlOoI
;
reg
CORETSE_AHBoOoI
;
reg
CORETSE_AHBiOoI
;
reg
CORETSE_AHBOIoI
;
wire
CORETSE_AHBIIoI
;
wire
CORETSE_AHBlIoI
;
wire
CORETSE_AHBoIoI
;
reg
CORETSE_AHBolOI
;
wire
[
RABITS
:
0
]
CORETSE_AHBilOI
;
reg
CORETSE_AHBiIoI
;
//      generated as part of synthesis results.
wire
[
(
RABITS
-
1
)
:
0
]
#
1000
CORETSE_AHBI0i
=
(
{
RABITS
{
~
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBlIoI
)
}
}
&
CORETSE_AHBOI1I
[
(
RABITS
+
1
)
:
CORETSE_AHBlo1
]
)
|
(
{
RABITS
{
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBlIoI
)
}
}
&
CORETSE_AHBiIII
[
(
RABITS
-
1
)
:
0
]
)
;
wire
#
1000
CORETSE_AHBO0i
=
~
(
CORETSE_AHBOl1I
&
~
CORETSE_AHBO01I
)
|
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBlIoI
)
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
1
]
<=
#
1000
1
'b
0
;
else
if
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBIIoI
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
1
]
<=
#
1000
CORETSE_AHBIlII
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
1
]
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
(
CORETSE_AHBiO1I
[
CORETSE_AHBlo1
-
1
:
0
]
==
{
CORETSE_AHBlo1
{
1
'h
0
}
}
)
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
1
]
<=
#
1000
CORETSE_AHBO1o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
]
<=
#
1000
1
'b
0
;
else
if
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBIIoI
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
]
<=
#
1000
CORETSE_AHBIlII
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
]
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
CORETSE_AHBO1o
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
]
<=
#
1000
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
CORETSE_AHBI1o
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
]
<=
#
1000
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+:
CORETSE_AHBlo1
]
<=
#
1000
{
CORETSE_AHBlo1
{
1
'h
0
}
}
;
else
if
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBIIoI
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+:
CORETSE_AHBlo1
]
<=
#
1000
CORETSE_AHBIlII
[
CORETSE_AHBIo1
+:
CORETSE_AHBlo1
]
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
CORETSE_AHBO1o
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+:
CORETSE_AHBlo1
]
<=
#
1000
{
CORETSE_AHBlo1
{
1
'h
0
}
}
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
CORETSE_AHBI1o
)
CORETSE_AHBl0i
[
CORETSE_AHBIo1
+:
CORETSE_AHBlo1
]
<=
#
1000
(
(
CORETSE_AHBIo1
/
8
)
-
1
)
-
CORETSE_AHBiO1I
[
(
CORETSE_AHBlo1
-
1
)
:
0
]
;
end
generate
genvar
CORETSE_AHBOloI
;
for
(
CORETSE_AHBOloI
=
0
;
CORETSE_AHBOloI
<
(
CORETSE_AHBIo1
/
8
)
;
CORETSE_AHBOloI
=
CORETSE_AHBOloI
+
1
)
begin
:
CORETSE_AHBIloI
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl0i
[
8
*
(
CORETSE_AHBOloI
+
1
)
-
1
:
CORETSE_AHBOloI
*
8
]
<=
#
1000
{
8
{
1
'h
0
}
}
;
else
if
(
~
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBIIoI
)
CORETSE_AHBl0i
[
8
*
(
CORETSE_AHBOloI
+
1
)
-
1
:
CORETSE_AHBOloI
*
8
]
<=
#
1000
CORETSE_AHBIlII
[
8
*
(
CORETSE_AHBOloI
+
1
)
-
1
:
CORETSE_AHBOloI
*
8
]
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
CORETSE_AHBiO1I
[
CORETSE_AHBlo1
-
1
:
0
]
==
CORETSE_AHBOloI
)
CORETSE_AHBl0i
[
8
*
(
CORETSE_AHBOloI
+
1
)
-
1
:
CORETSE_AHBOloI
*
8
]
<=
#
1000
CORETSE_AHBo0o
;
end
end
endgenerate
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBiI1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
(
CORETSE_AHBI1o
|
CORETSE_AHBO01I
)
&
CORETSE_AHBi0o
)
CORETSE_AHBiI1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBO1o
)
CORETSE_AHBiI1I
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
assign
CORETSE_AHBoI1I
=
(
CORETSE_AHBiI1I
|
CORETSE_AHBO1o
)
&
~
CORETSE_AHBO01I
&
CORETSE_AHBi0o
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOl1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBOl1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI1I
;
end
assign
CORETSE_AHBO01I
=
(
CORETSE_AHBOI1I
[
(
RABITS
+
CORETSE_AHBlo1
)
-
1
:
CORETSE_AHBlo1
]
==
CORETSE_AHBi01I
[
(
RABITS
-
1
)
:
0
]
)
&
(
CORETSE_AHBOI1I
[
RABITS
+
CORETSE_AHBlo1
]
!=
CORETSE_AHBi01I
[
RABITS
]
)
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBI01I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBI01I
<=
#
CORETSE_AHBIoII
CORETSE_AHBO01I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBO01I
)
CORETSE_AHBoIOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBo01I
)
CORETSE_AHBoIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
assign
CORETSE_AHBIl1I
=
CORETSE_AHBOI1I
+
1
'b
1
;
assign
CORETSE_AHBll1I
=
{
CORETSE_AHBOI1I
[
(
RABITS
+
CORETSE_AHBlo1
)
:
CORETSE_AHBlo1
]
,
{
CORETSE_AHBlo1
{
1
'h
0
}
}
}
+
(
CORETSE_AHBIo1
/
8
)
;
assign
CORETSE_AHBiO1I
=
(
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBoIoI
)
?
{
CORETSE_AHBiIII
[
RABITS
:
0
]
,
{
CORETSE_AHBlo1
{
1
'h
0
}
}
}
:
(
CORETSE_AHBol1I
)
?
CORETSE_AHBII1I
:
(
CORETSE_AHBO01I
)
?
CORETSE_AHBOI1I
:
(
CORETSE_AHBOl1I
&
CORETSE_AHBlI1I
)
?
CORETSE_AHBll1I
:
(
CORETSE_AHBoI1I
&
~
CORETSE_AHBO1o
)
?
CORETSE_AHBIl1I
:
CORETSE_AHBOI1I
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOI1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBOI1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBlI1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBlI1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1o
;
end
generate
if
(
CORETSE_AHBoOI
==
1
)
begin
assign
CORETSE_AHBlloI
=
CORETSE_AHBoo1I
;
end
endgenerate
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBi01I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoO1I
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBOo1I
&
~
CORETSE_AHBoii
)
CORETSE_AHBi01I
<=
#
CORETSE_AHBIoII
CORETSE_AHBioi
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBII1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBO1o
&
~
CORETSE_AHBol1I
)
CORETSE_AHBII1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBol1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
(
CORETSE_AHBoo1I
|
(
~
CORETSE_AHBIIOI
&
(
CORETSE_AHBOl1I
&
CORETSE_AHBoI1I
)
)
|
(
CORETSE_AHBO01I
&
(
CORETSE_AHBOl1I
|
CORETSE_AHBoI1I
)
)
)
)
CORETSE_AHBol1I
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBO1o
&
~
CORETSE_AHBO01I
)
CORETSE_AHBol1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBiIoI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiIoI
<=
(
CORETSE_AHBi1o
&
CORETSE_AHBo1o
)
|
(
CORETSE_AHBiIoI
&
!
CORETSE_AHBii1I
)
;
end
assign
CORETSE_AHBOOoI
=
(
CORETSE_AHBo1o
&
~
CORETSE_AHBli1I
)
|
(
CORETSE_AHBoi1I
&
CORETSE_AHBii1I
)
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBli1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBli1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoi1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBoi1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBli1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBii1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBii1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1o
;
end
assign
CORETSE_AHBlOoI
=
CORETSE_AHBOOoI
&
(
(
|
(
(
{
CORETSE_AHBiIoI
,
CORETSE_AHBl1o
[
32
:
16
]
}
~^
CORETSE_AHBOoOI
)
&
~
CORETSE_AHBIoOI
)
)
|
(
(
CORETSE_AHBl1o
[
15
:
0
]
<
16
'd
64
)
&
CORETSE_AHBloOI
)
|
CORETSE_AHBOoo
)
;
assign
CORETSE_AHBio1I
=
CORETSE_AHBOOoI
&
~
CORETSE_AHBlOoI
;
assign
CORETSE_AHBoo1I
=
CORETSE_AHBlOoI
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIi1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO1I
;
else
if
(
CORETSE_AHBl0o
&
~
CORETSE_AHBOi1I
)
CORETSE_AHBIi1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO1I
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoI1I
&
~
(
&
CORETSE_AHBIi1I
)
)
CORETSE_AHBIi1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi1I
+
1
;
end
assign
CORETSE_AHBIOoI
=
(
CORETSE_AHBiIII
[
RABITS
+
1
]
&
CORETSE_AHBlIoI
)
|
(
CORETSE_AHBio1I
&
~
CORETSE_AHBI01I
)
|
(
(
CORETSE_AHBIi1I
[
(
RABITS
+
CORETSE_AHBlo1
)
-
1
:
CORETSE_AHBlo1
]
>=
CORETSE_AHBi1OI
)
&
~
(
&
CORETSE_AHBi1OI
)
&
(
&
CORETSE_AHBiO1I
[
CORETSE_AHBlo1
-
1
:
0
]
)
&
~
CORETSE_AHBI01I
)
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBil1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBoO1I
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBIOoI
)
CORETSE_AHBil1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO1I
[
(
RABITS
+
CORETSE_AHBlo1
)
:
CORETSE_AHBlo1
]
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBlii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBI11I
)
CORETSE_AHBlii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBlii
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIii
<=
#
CORETSE_AHBIoII
CORETSE_AHBoO1I
;
else
if
(
CORETSE_AHBl0o
&
~
CORETSE_AHBI11I
&
~
CORETSE_AHBlii
)
CORETSE_AHBIii
<=
#
CORETSE_AHBIoII
CORETSE_AHBil1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBo11I
)
CORETSE_AHBIOOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBIOOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBiii
<=
#
CORETSE_AHBIoII
CORETSE_AHBoO1I
;
else
if
(
CORETSE_AHBl0o
&
~
CORETSE_AHBo11I
&
~
CORETSE_AHBIOOI
)
CORETSE_AHBiii
<=
#
CORETSE_AHBIoII
CORETSE_AHBil1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoO1I
;
else
if
(
CORETSE_AHBl0o
&
~
CORETSE_AHBo11I
&
~
CORETSE_AHBIOOI
)
CORETSE_AHBOOOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi01I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
~
CORETSE_AHBOo1I
)
CORETSE_AHBoii
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBOo1I
)
CORETSE_AHBoii
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBO1o
&
CORETSE_AHBlo1I
)
CORETSE_AHBIIOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBl0o
&
(
CORETSE_AHBI1o
|
~
CORETSE_AHBOi1I
)
&
~
CORETSE_AHBlo1I
)
CORETSE_AHBIIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOi1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBO1o
&
CORETSE_AHBlo1I
)
CORETSE_AHBOi1I
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBI1o
)
CORETSE_AHBOi1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl01I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl01I
<=
#
CORETSE_AHBIoII
CORETSE_AHBooOI
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBo01I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo01I
<=
#
CORETSE_AHBIoII
CORETSE_AHBl01I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBO11I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO11I
<=
#
CORETSE_AHBIoII
CORETSE_AHBooi
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBI11I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI11I
<=
#
CORETSE_AHBIoII
CORETSE_AHBO11I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl11I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl11I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOOI
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBo11I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo11I
<=
#
CORETSE_AHBIoII
CORETSE_AHBl11I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBi11I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi11I
<=
#
CORETSE_AHBIoII
CORETSE_AHBOii
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOo1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOo1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi11I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIo1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIo1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBlOII
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBlo1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlo1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoOoI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoOoI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOlII
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBiOoI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiOoI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOoI
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOIoI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOIoI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOoI
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBolOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBolOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIoI
;
end
assign
CORETSE_AHBIIoI
=
CORETSE_AHBiOoI
&
~
CORETSE_AHBOIoI
;
assign
CORETSE_AHBlIoI
=
CORETSE_AHBOIoI
&
~
CORETSE_AHBolOI
;
assign
CORETSE_AHBoIoI
=
CORETSE_AHBlIoI
|
CORETSE_AHBIIoI
;
assign
CORETSE_AHBilOI
=
CORETSE_AHBOI1I
[
(
RABITS
+
CORETSE_AHBlo1
)
:
CORETSE_AHBlo1
]
;
endmodule
