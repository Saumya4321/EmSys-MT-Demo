// REVISION    : $Revision: 1.1 $
//              Mentor Proprietary and Confidential
//              Copyright (c) 2000, Mentor Intellectual Property Development
`timescale 1ns/1ns
module
pemstat_ladd
(
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
,
CORETSE_AHBi10i
,
CORETSE_AHBOo0i
,
CORETSE_AHBoIIi
,
CORETSE_AHBl1li
,
CORETSE_AHBiIIi
,
CORETSE_AHBlIIi
,
CORETSE_AHBIo0i
,
CORETSE_AHBoOIi
)
;
input
CORETSE_AHBi1Oi
,
CORETSE_AHBo1Oi
;
input
CORETSE_AHBi10i
;
input
[
15
:
0
]
CORETSE_AHBOo0i
;
input
CORETSE_AHBoIIi
;
input
[
30
:
0
]
CORETSE_AHBl1li
;
input
CORETSE_AHBiIIi
;
input
CORETSE_AHBlIIi
;
output
[
30
:
0
]
CORETSE_AHBIo0i
;
output
CORETSE_AHBoOIi
;
reg
CORETSE_AHBoOIi
;
parameter
CORETSE_AHBIoII
=
1
;
wire
[
24
:
0
]
CORETSE_AHBlo0i
;
reg
[
23
:
0
]
CORETSE_AHBoo0i
;
assign
CORETSE_AHBlo0i
[
24
:
0
]
=
CORETSE_AHBoo0i
[
23
:
0
]
+
{
8
'h
0
,
CORETSE_AHBOo0i
[
15
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBoo0i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
24
'h
0
;
else
if
(
CORETSE_AHBoIIi
)
CORETSE_AHBoo0i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1li
[
23
:
0
]
;
else
if
(
CORETSE_AHBi10i
&
CORETSE_AHBlIIi
)
CORETSE_AHBoo0i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
{
8
'h
0
,
CORETSE_AHBOo0i
[
15
:
0
]
}
;
else
if
(
CORETSE_AHBi10i
)
CORETSE_AHBoo0i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBlo0i
[
23
:
0
]
;
else
if
(
CORETSE_AHBlIIi
)
CORETSE_AHBoo0i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
24
'h
0
;
else
CORETSE_AHBoo0i
[
23
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0i
[
23
:
0
]
;
end
assign
CORETSE_AHBIo0i
[
30
:
0
]
=
{
7
'h
0
,
CORETSE_AHBoo0i
[
23
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo1Oi
or
posedge
CORETSE_AHBi1Oi
)
begin
if
(
CORETSE_AHBi1Oi
)
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBiIIi
)
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi10i
&
CORETSE_AHBlo0i
[
24
]
)
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
CORETSE_AHBoOIi
<=
#
CORETSE_AHBIoII
CORETSE_AHBoOIi
;
end
endmodule
