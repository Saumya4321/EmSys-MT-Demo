// REVISION    : $Revision: 1.10 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxfif
#
(
parameter
TABITS
=
12
,
parameter
RABITS
=
12
,
parameter
CORETSE_AHBIo1
=
32
,
parameter
CORETSE_AHBlo1
=
$clog2
(
CORETSE_AHBIo1
/
8
)
,
parameter
CORETSE_AHBoOI
=
0
)
(
CORETSE_AHBIi0
,
CORETSE_AHBoo1
,
CORETSE_AHBio1
,
CORETSE_AHBOi1
,
CORETSE_AHBIi1
,
CORETSE_AHBli1
,
CORETSE_AHBoi1
,
CORETSE_AHBii1
,
CORETSE_AHBOOo
,
CORETSE_AHBIOo
,
CORETSE_AHBlOo
,
CORETSE_AHBoOo
,
CORETSE_AHBiOo
,
CORETSE_AHBOIo
,
CORETSE_AHBIIo
,
CORETSE_AHBlIo
,
CORETSE_AHBoIo
,
CORETSE_AHBiIo
,
CORETSE_AHBOlo
,
CORETSE_AHBIlo
,
CORETSE_AHBoi0
,
CORETSE_AHBllo
,
CORETSE_AHBolo
,
CORETSE_AHBilo
,
CORETSE_AHBO0o
,
CORETSE_AHBI0o
,
CORETSE_AHBii0
,
CORETSE_AHBl0o
,
CORETSE_AHBo0o
,
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
,
CORETSE_AHBl1o
,
CORETSE_AHBo1o
,
CORETSE_AHBi1o
,
CORETSE_AHBOoo
,
CORETSE_AHBIoo
,
CORETSE_AHBloo
,
CORETSE_AHBooo
,
CORETSE_AHBioo
,
CORETSE_AHBOio
,
CORETSE_AHBIio
,
CORETSE_AHBlio
,
CORETSE_AHBoio
,
CORETSE_AHBiio
,
CORETSE_AHBOOi
,
CORETSE_AHBIOi
,
CORETSE_AHBlOi
,
CORETSE_AHBoOi
,
CORETSE_AHBiOi
,
CORETSE_AHBOIi
,
CORETSE_AHBIIi
,
CORETSE_AHBlIi
,
CORETSE_AHBoIi
,
CORETSE_AHBiIi
,
CORETSE_AHBOli
,
CORETSE_AHBIli
,
CORETSE_AHBlli
,
CORETSE_AHBoli
,
CORETSE_AHBili
,
CORETSE_AHBO0i
,
CORETSE_AHBI0i
,
CORETSE_AHBl0i
,
CORETSE_AHBo0i
,
CORETSE_AHBi0i
,
CORETSE_AHBO1i
,
CORETSE_AHBI1i
)
;
input
CORETSE_AHBIi0
;
input
CORETSE_AHBoo1
;
input
CORETSE_AHBio1
;
input
CORETSE_AHBOi1
;
input
CORETSE_AHBIi1
;
input
CORETSE_AHBli1
;
input
[
7
:
0
]
CORETSE_AHBoi1
;
input
[
31
:
0
]
CORETSE_AHBii1
;
input
CORETSE_AHBOOo
;
input
[
(
CORETSE_AHBIo1
-
1
)
:
0
]
CORETSE_AHBIOo
;
input
CORETSE_AHBlOo
;
input
CORETSE_AHBoOo
;
input
[
1
:
0
]
CORETSE_AHBiOo
;
input
CORETSE_AHBOIo
;
input
CORETSE_AHBIIo
;
input
[
1
:
0
]
CORETSE_AHBlIo
;
input
CORETSE_AHBoIo
;
input
CORETSE_AHBiIo
;
input
CORETSE_AHBOlo
;
input
CORETSE_AHBIlo
;
input
CORETSE_AHBoi0
;
input
CORETSE_AHBllo
;
input
CORETSE_AHBolo
;
input
CORETSE_AHBilo
;
input
CORETSE_AHBO0o
;
input
CORETSE_AHBI0o
;
input
CORETSE_AHBii0
;
input
CORETSE_AHBl0o
;
input
[
7
:
0
]
CORETSE_AHBo0o
;
input
CORETSE_AHBi0o
;
input
CORETSE_AHBO1o
;
input
CORETSE_AHBI1o
;
input
[
32
:
0
]
CORETSE_AHBl1o
;
input
CORETSE_AHBo1o
;
input
CORETSE_AHBi1o
;
input
CORETSE_AHBOoo
;
input
CORETSE_AHBIoo
;
output
CORETSE_AHBloo
;
output
CORETSE_AHBooo
;
output
[
(
CORETSE_AHBIo1
-
1
)
:
0
]
CORETSE_AHBioo
;
output
CORETSE_AHBOio
;
output
CORETSE_AHBIio
;
output
[
1
:
0
]
CORETSE_AHBlio
;
output
CORETSE_AHBoio
;
output
[
7
:
0
]
CORETSE_AHBiio
;
output
CORETSE_AHBOOi
;
output
CORETSE_AHBIOi
;
output
CORETSE_AHBlOi
;
output
CORETSE_AHBoOi
;
output
CORETSE_AHBiOi
;
output
CORETSE_AHBOIi
;
output
CORETSE_AHBIIi
;
output
CORETSE_AHBlIi
;
output
CORETSE_AHBoIi
;
output
CORETSE_AHBiIi
;
output
CORETSE_AHBOli
;
output
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBIli
;
output
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBlli
;
output
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBoli
;
input
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBili
;
output
CORETSE_AHBO0i
;
output
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBI0i
;
output
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBl0i
;
output
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBo0i
;
input
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBi0i
;
output
[
31
:
0
]
CORETSE_AHBO1i
;
output
CORETSE_AHBI1i
;
wire
CORETSE_AHBl1i
;
wire
[
TABITS
:
0
]
CORETSE_AHBo1i
;
wire
CORETSE_AHBi1i
;
wire
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBIli
;
wire
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBlli
;
wire
CORETSE_AHBOli
;
wire
[
TABITS
:
0
]
CORETSE_AHBOoi
;
wire
CORETSE_AHBIoi
;
wire
CORETSE_AHBloi
;
wire
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBili
;
wire
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBoli
;
wire
CORETSE_AHBooi
;
wire
[
RABITS
:
0
]
CORETSE_AHBioi
;
wire
CORETSE_AHBOii
;
wire
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBI0i
;
wire
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBl0i
;
wire
CORETSE_AHBO0i
;
wire
[
RABITS
:
0
]
CORETSE_AHBIii
;
wire
CORETSE_AHBlii
;
wire
CORETSE_AHBoii
;
wire
[
(
CORETSE_AHBIo1
+
4
)
-
1
:
0
]
CORETSE_AHBi0i
;
wire
[
(
RABITS
-
1
)
:
0
]
CORETSE_AHBo0i
;
wire
[
RABITS
:
0
]
CORETSE_AHBiii
;
wire
[
RABITS
:
0
]
CORETSE_AHBOOOI
;
wire
CORETSE_AHBIOOI
;
wire
CORETSE_AHBlOOI
;
wire
CORETSE_AHBoOOI
;
wire
CORETSE_AHBiOOI
;
wire
CORETSE_AHBOIOI
;
wire
CORETSE_AHBIIOI
;
wire
CORETSE_AHBlIOI
;
wire
CORETSE_AHBoIOI
;
wire
CORETSE_AHBiIOI
;
wire
[
TABITS
:
0
]
CORETSE_AHBOlOI
;
wire
CORETSE_AHBIlOI
;
wire
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBllOI
;
wire
CORETSE_AHBolOI
;
wire
[
RABITS
:
0
]
CORETSE_AHBilOI
;
wire
CORETSE_AHBO0OI
;
wire
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBI0OI
;
wire
[
15
:
0
]
CORETSE_AHBl0OI
;
wire
[
RABITS
:
0
]
CORETSE_AHBo0OI
;
wire
[
RABITS
:
0
]
CORETSE_AHBi0OI
;
wire
CORETSE_AHBO1OI
;
wire
CORETSE_AHBI1OI
;
wire
[
TABITS
:
0
]
CORETSE_AHBl1OI
;
wire
[
TABITS
:
0
]
CORETSE_AHBo1OI
;
wire
[
RABITS
-
1
:
0
]
CORETSE_AHBi1OI
;
wire
[
17
:
0
]
CORETSE_AHBOoOI
;
wire
[
17
:
0
]
CORETSE_AHBIoOI
;
wire
CORETSE_AHBloOI
;
wire
CORETSE_AHBooOI
;
wire
CORETSE_AHBioOI
;
wire
CORETSE_AHBOiOI
;
wire
CORETSE_AHBIiOI
;
wire
CORETSE_AHBliOI
;
wire
CORETSE_AHBoiOI
;
wire
CORETSE_AHBiiOI
;
wire
CORETSE_AHBOOII
;
wire
CORETSE_AHBIOII
;
wire
CORETSE_AHBlOII
;
wire
CORETSE_AHBoOII
;
wire
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBiOII
;
wire
CORETSE_AHBOIII
;
wire
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIIII
;
wire
[
(
TABITS
+
1
)
:
0
]
CORETSE_AHBlIII
;
wire
CORETSE_AHBoIII
;
wire
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBiIII
;
wire
CORETSE_AHBOlII
;
wire
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBIlII
;
wire
[
(
RABITS
+
1
)
:
0
]
CORETSE_AHBllII
;
wire
CORETSE_AHBolII
;
wire
[
31
:
0
]
CORETSE_AHBO1i
;
wire
CORETSE_AHBI1i
;
wire
CORETSE_AHBilII
;
wire
CORETSE_AHBO0II
;
wire
CORETSE_AHBI0II
;
wire
CORETSE_AHBl0II
;
wire
CORETSE_AHBo0II
;
amcxtfif_fab
#
(
.TABITS
(
TABITS
)
,
.CORETSE_AHBIo1
(
CORETSE_AHBIo1
)
,
.CORETSE_AHBlo1
(
CORETSE_AHBlo1
)
)
CORETSE_AHBi0II
(
.CORETSE_AHBOOo
(
CORETSE_AHBOOo
)
,
.CORETSE_AHBilII
(
CORETSE_AHBilII
)
,
.CORETSE_AHBiiOI
(
CORETSE_AHBiiOI
)
,
.CORETSE_AHBIOo
(
CORETSE_AHBIOo
)
,
.CORETSE_AHBlOo
(
CORETSE_AHBlOo
)
,
.CORETSE_AHBoOo
(
CORETSE_AHBoOo
)
,
.CORETSE_AHBiOo
(
CORETSE_AHBiOo
)
,
.CORETSE_AHBOIo
(
CORETSE_AHBOIo
)
,
.CORETSE_AHBIIo
(
CORETSE_AHBIIo
)
,
.CORETSE_AHBlIo
(
CORETSE_AHBlIo
)
,
.CORETSE_AHBoIo
(
CORETSE_AHBoIo
)
,
.CORETSE_AHBiIo
(
CORETSE_AHBiIo
)
,
.CORETSE_AHBl1i
(
CORETSE_AHBl1i
)
,
.CORETSE_AHBo1i
(
CORETSE_AHBo1i
)
,
.CORETSE_AHBi1i
(
CORETSE_AHBi1i
)
,
.CORETSE_AHBl1OI
(
CORETSE_AHBl1OI
)
,
.CORETSE_AHBo1OI
(
CORETSE_AHBo1OI
)
,
.CORETSE_AHBiOII
(
CORETSE_AHBiOII
)
,
.CORETSE_AHBOIII
(
CORETSE_AHBOIII
)
,
.CORETSE_AHBIIII
(
CORETSE_AHBIIII
)
,
.CORETSE_AHBoOOI
(
CORETSE_AHBoOOI
)
,
.CORETSE_AHBIli
(
CORETSE_AHBIli
)
,
.CORETSE_AHBlli
(
CORETSE_AHBlli
)
,
.CORETSE_AHBOli
(
CORETSE_AHBOli
)
,
.CORETSE_AHBloo
(
CORETSE_AHBloo
)
,
.CORETSE_AHBooo
(
CORETSE_AHBooo
)
,
.CORETSE_AHBOoi
(
CORETSE_AHBOoi
)
,
.CORETSE_AHBIoi
(
CORETSE_AHBIoi
)
,
.CORETSE_AHBloi
(
CORETSE_AHBloi
)
,
.CORETSE_AHBiIOI
(
CORETSE_AHBiIOI
)
,
.CORETSE_AHBOlOI
(
CORETSE_AHBOlOI
)
)
;
amcxtfif_sys
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
,
.TABITS
(
TABITS
)
,
.CORETSE_AHBIo1
(
CORETSE_AHBIo1
)
,
.CORETSE_AHBlo1
(
CORETSE_AHBlo1
)
)
CORETSE_AHBO1II
(
.CORETSE_AHBoi0
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBllo
(
CORETSE_AHBllo
)
,
.CORETSE_AHBO0II
(
CORETSE_AHBO0II
)
,
.CORETSE_AHBOOII
(
CORETSE_AHBOOII
)
,
.CORETSE_AHBili
(
CORETSE_AHBili
)
,
.CORETSE_AHBolo
(
CORETSE_AHBolo
)
,
.CORETSE_AHBilo
(
CORETSE_AHBilo
)
,
.CORETSE_AHBO0o
(
CORETSE_AHBO0o
)
,
.CORETSE_AHBI0o
(
CORETSE_AHBI0o
)
,
.CORETSE_AHBOoi
(
CORETSE_AHBOoi
)
,
.CORETSE_AHBIoi
(
CORETSE_AHBIoi
)
,
.CORETSE_AHBloi
(
CORETSE_AHBloi
)
,
.CORETSE_AHBlIII
(
CORETSE_AHBlIII
)
,
.CORETSE_AHBoIII
(
CORETSE_AHBoIII
)
,
.CORETSE_AHBiOOI
(
CORETSE_AHBiOOI
)
,
.CORETSE_AHBoli
(
CORETSE_AHBoli
)
,
.CORETSE_AHBiio
(
CORETSE_AHBiio
)
,
.CORETSE_AHBOOi
(
CORETSE_AHBOOi
)
,
.CORETSE_AHBIOi
(
CORETSE_AHBIOi
)
,
.CORETSE_AHBlOi
(
CORETSE_AHBlOi
)
,
.CORETSE_AHBoOi
(
CORETSE_AHBoOi
)
,
.CORETSE_AHBiOi
(
CORETSE_AHBiOi
)
,
.CORETSE_AHBOIi
(
CORETSE_AHBOIi
)
,
.CORETSE_AHBIIi
(
CORETSE_AHBIIi
)
,
.CORETSE_AHBl1i
(
CORETSE_AHBl1i
)
,
.CORETSE_AHBo1i
(
CORETSE_AHBo1i
)
,
.CORETSE_AHBi1i
(
CORETSE_AHBi1i
)
,
.CORETSE_AHBIlOI
(
CORETSE_AHBIlOI
)
,
.CORETSE_AHBllOI
(
CORETSE_AHBllOI
)
)
;
amcxrfif_fab
#
(
.RABITS
(
RABITS
)
,
.CORETSE_AHBIo1
(
CORETSE_AHBIo1
)
,
.CORETSE_AHBlo1
(
CORETSE_AHBlo1
)
)
CORETSE_AHBI1II
(
.CORETSE_AHBOlo
(
CORETSE_AHBOlo
)
,
.CORETSE_AHBI0II
(
CORETSE_AHBI0II
)
,
.CORETSE_AHBIOII
(
CORETSE_AHBIOII
)
,
.CORETSE_AHBIlo
(
CORETSE_AHBIlo
)
,
.CORETSE_AHBi0i
(
CORETSE_AHBi0i
)
,
.CORETSE_AHBIii
(
CORETSE_AHBIii
)
,
.CORETSE_AHBlii
(
CORETSE_AHBlii
)
,
.CORETSE_AHBoii
(
CORETSE_AHBoii
)
,
.CORETSE_AHBllII
(
CORETSE_AHBllII
)
,
.CORETSE_AHBolII
(
CORETSE_AHBolII
)
,
.CORETSE_AHBOIOI
(
CORETSE_AHBOIOI
)
,
.CORETSE_AHBo0i
(
CORETSE_AHBo0i
)
,
.CORETSE_AHBioo
(
CORETSE_AHBioo
)
,
.CORETSE_AHBOio
(
CORETSE_AHBOio
)
,
.CORETSE_AHBIio
(
CORETSE_AHBIio
)
,
.CORETSE_AHBlio
(
CORETSE_AHBlio
)
,
.CORETSE_AHBoio
(
CORETSE_AHBoio
)
,
.CORETSE_AHBooi
(
CORETSE_AHBooi
)
,
.CORETSE_AHBioi
(
CORETSE_AHBioi
)
,
.CORETSE_AHBOii
(
CORETSE_AHBOii
)
,
.CORETSE_AHBO0OI
(
CORETSE_AHBO0OI
)
,
.CORETSE_AHBI0OI
(
CORETSE_AHBI0OI
)
)
;
amcxrfif_sys
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
,
.RABITS
(
RABITS
)
,
.CORETSE_AHBIo1
(
CORETSE_AHBIo1
)
,
.CORETSE_AHBlo1
(
CORETSE_AHBlo1
)
)
CORETSE_AHBl1II
(
.CORETSE_AHBii0
(
CORETSE_AHBii0
)
,
.CORETSE_AHBl0o
(
CORETSE_AHBl0o
)
,
.CORETSE_AHBl0II
(
CORETSE_AHBl0II
)
,
.CORETSE_AHBlOII
(
CORETSE_AHBlOII
)
,
.CORETSE_AHBi1OI
(
CORETSE_AHBi1OI
)
,
.CORETSE_AHBOoOI
(
CORETSE_AHBOoOI
)
,
.CORETSE_AHBIoOI
(
CORETSE_AHBIoOI
)
,
.CORETSE_AHBloOI
(
CORETSE_AHBloOI
)
,
.CORETSE_AHBooOI
(
CORETSE_AHBooOI
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBo0o
)
,
.CORETSE_AHBi0o
(
CORETSE_AHBi0o
)
,
.CORETSE_AHBO1o
(
CORETSE_AHBO1o
)
,
.CORETSE_AHBI1o
(
CORETSE_AHBI1o
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBi1o
(
CORETSE_AHBi1o
)
,
.CORETSE_AHBOoo
(
CORETSE_AHBOoo
)
,
.CORETSE_AHBooi
(
CORETSE_AHBooi
)
,
.CORETSE_AHBlOOI
(
CORETSE_AHBlOOI
)
,
.CORETSE_AHBioi
(
CORETSE_AHBioi
)
,
.CORETSE_AHBOii
(
CORETSE_AHBOii
)
,
.CORETSE_AHBiIII
(
CORETSE_AHBiIII
)
,
.CORETSE_AHBOlII
(
CORETSE_AHBOlII
)
,
.CORETSE_AHBIlII
(
CORETSE_AHBIlII
)
,
.CORETSE_AHBIIOI
(
CORETSE_AHBIIOI
)
,
.CORETSE_AHBoIOI
(
CORETSE_AHBoIOI
)
,
.CORETSE_AHBI0i
(
CORETSE_AHBI0i
)
,
.CORETSE_AHBl0i
(
CORETSE_AHBl0i
)
,
.CORETSE_AHBO0i
(
CORETSE_AHBO0i
)
,
.CORETSE_AHBIii
(
CORETSE_AHBIii
)
,
.CORETSE_AHBlii
(
CORETSE_AHBlii
)
,
.CORETSE_AHBiii
(
CORETSE_AHBiii
)
,
.CORETSE_AHBOOOI
(
CORETSE_AHBOOOI
)
,
.CORETSE_AHBIOOI
(
CORETSE_AHBIOOI
)
,
.CORETSE_AHBoii
(
CORETSE_AHBoii
)
,
.CORETSE_AHBolOI
(
CORETSE_AHBolOI
)
,
.CORETSE_AHBilOI
(
CORETSE_AHBilOI
)
)
;
amcxtfif_wtm
#
(
.RABITS
(
RABITS
)
)
CORETSE_AHBo1II
(
.CORETSE_AHBoi0
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBllo
(
CORETSE_AHBllo
)
,
.CORETSE_AHBo0II
(
CORETSE_AHBo0II
)
,
.CORETSE_AHBoOII
(
CORETSE_AHBoOII
)
,
.CORETSE_AHBl0OI
(
CORETSE_AHBl0OI
)
,
.CORETSE_AHBo0OI
(
CORETSE_AHBo0OI
)
,
.CORETSE_AHBi0OI
(
CORETSE_AHBi0OI
)
,
.CORETSE_AHBO1OI
(
CORETSE_AHBO1OI
)
,
.CORETSE_AHBI1OI
(
CORETSE_AHBI1OI
)
,
.CORETSE_AHBIoo
(
CORETSE_AHBIoo
)
,
.CORETSE_AHBiii
(
CORETSE_AHBiii
)
,
.CORETSE_AHBOOOI
(
CORETSE_AHBOOOI
)
,
.CORETSE_AHBIOOI
(
CORETSE_AHBIOOI
)
,
.CORETSE_AHBlIOI
(
CORETSE_AHBlIOI
)
,
.CORETSE_AHBlIi
(
CORETSE_AHBlIi
)
,
.CORETSE_AHBoIi
(
CORETSE_AHBoIi
)
,
.CORETSE_AHBiIi
(
CORETSE_AHBiIi
)
,
.CORETSE_AHBlOOI
(
CORETSE_AHBlOOI
)
)
;
amcxfif_hst
#
(
.TABITS
(
TABITS
)
,
.RABITS
(
RABITS
)
,
.CORETSE_AHBIo1
(
CORETSE_AHBIo1
)
,
.CORETSE_AHBlo1
(
CORETSE_AHBlo1
)
)
CORETSE_AHBi1II
(
.CORETSE_AHBio1
(
CORETSE_AHBio1
)
,
.CORETSE_AHBOi1
(
CORETSE_AHBOi1
)
,
.CORETSE_AHBIi1
(
CORETSE_AHBIi1
)
,
.CORETSE_AHBli1
(
CORETSE_AHBli1
)
,
.CORETSE_AHBoi1
(
CORETSE_AHBoi1
)
,
.CORETSE_AHBii1
(
CORETSE_AHBii1
)
,
.CORETSE_AHBoOOI
(
CORETSE_AHBoOOI
)
,
.CORETSE_AHBiOOI
(
CORETSE_AHBiOOI
)
,
.CORETSE_AHBOIOI
(
CORETSE_AHBOIOI
)
,
.CORETSE_AHBIIOI
(
CORETSE_AHBIIOI
)
,
.CORETSE_AHBlIOI
(
CORETSE_AHBlIOI
)
,
.CORETSE_AHBoIOI
(
CORETSE_AHBoIOI
)
,
.CORETSE_AHBiIOI
(
CORETSE_AHBiIOI
)
,
.CORETSE_AHBOlOI
(
CORETSE_AHBOlOI
)
,
.CORETSE_AHBIlOI
(
CORETSE_AHBIlOI
)
,
.CORETSE_AHBllOI
(
CORETSE_AHBllOI
)
,
.CORETSE_AHBolOI
(
CORETSE_AHBolOI
)
,
.CORETSE_AHBilOI
(
CORETSE_AHBilOI
)
,
.CORETSE_AHBO0OI
(
CORETSE_AHBO0OI
)
,
.CORETSE_AHBI0OI
(
CORETSE_AHBI0OI
)
,
.CORETSE_AHBl1OI
(
CORETSE_AHBl1OI
)
,
.CORETSE_AHBo1OI
(
CORETSE_AHBo1OI
)
,
.CORETSE_AHBi1OI
(
CORETSE_AHBi1OI
)
,
.CORETSE_AHBl0OI
(
CORETSE_AHBl0OI
)
,
.CORETSE_AHBo0OI
(
CORETSE_AHBo0OI
)
,
.CORETSE_AHBi0OI
(
CORETSE_AHBi0OI
)
,
.CORETSE_AHBO1OI
(
CORETSE_AHBO1OI
)
,
.CORETSE_AHBI1OI
(
CORETSE_AHBI1OI
)
,
.CORETSE_AHBOoOI
(
CORETSE_AHBOoOI
)
,
.CORETSE_AHBIoOI
(
CORETSE_AHBIoOI
)
,
.CORETSE_AHBloOI
(
CORETSE_AHBloOI
)
,
.CORETSE_AHBooOI
(
CORETSE_AHBooOI
)
,
.CORETSE_AHBioOI
(
CORETSE_AHBioOI
)
,
.CORETSE_AHBOiOI
(
CORETSE_AHBOiOI
)
,
.CORETSE_AHBIiOI
(
CORETSE_AHBIiOI
)
,
.CORETSE_AHBliOI
(
CORETSE_AHBliOI
)
,
.CORETSE_AHBoiOI
(
CORETSE_AHBoiOI
)
,
.CORETSE_AHBiiOI
(
CORETSE_AHBiiOI
)
,
.CORETSE_AHBOOII
(
CORETSE_AHBOOII
)
,
.CORETSE_AHBIOII
(
CORETSE_AHBIOII
)
,
.CORETSE_AHBlOII
(
CORETSE_AHBlOII
)
,
.CORETSE_AHBoOII
(
CORETSE_AHBoOII
)
,
.CORETSE_AHBiOII
(
CORETSE_AHBiOII
)
,
.CORETSE_AHBOIII
(
CORETSE_AHBOIII
)
,
.CORETSE_AHBIIII
(
CORETSE_AHBIIII
)
,
.CORETSE_AHBlIII
(
CORETSE_AHBlIII
)
,
.CORETSE_AHBoIII
(
CORETSE_AHBoIII
)
,
.CORETSE_AHBiIII
(
CORETSE_AHBiIII
)
,
.CORETSE_AHBOlII
(
CORETSE_AHBOlII
)
,
.CORETSE_AHBIlII
(
CORETSE_AHBIlII
)
,
.CORETSE_AHBllII
(
CORETSE_AHBllII
)
,
.CORETSE_AHBolII
(
CORETSE_AHBolII
)
,
.CORETSE_AHBO1i
(
CORETSE_AHBO1i
)
,
.CORETSE_AHBI1i
(
CORETSE_AHBI1i
)
)
;
amcxfif_clkrst
CORETSE_AHBOoII
(
.CORETSE_AHBIi0
(
CORETSE_AHBIi0
)
,
.CORETSE_AHBoo1
(
CORETSE_AHBoo1
)
,
.CORETSE_AHBoi0
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBii0
(
CORETSE_AHBii0
)
,
.CORETSE_AHBOOo
(
CORETSE_AHBOOo
)
,
.CORETSE_AHBOlo
(
CORETSE_AHBOlo
)
,
.CORETSE_AHBioOI
(
CORETSE_AHBioOI
)
,
.CORETSE_AHBOiOI
(
CORETSE_AHBOiOI
)
,
.CORETSE_AHBIiOI
(
CORETSE_AHBIiOI
)
,
.CORETSE_AHBliOI
(
CORETSE_AHBliOI
)
,
.CORETSE_AHBoiOI
(
CORETSE_AHBoiOI
)
,
.CORETSE_AHBilII
(
CORETSE_AHBilII
)
,
.CORETSE_AHBO0II
(
CORETSE_AHBO0II
)
,
.CORETSE_AHBI0II
(
CORETSE_AHBI0II
)
,
.CORETSE_AHBl0II
(
CORETSE_AHBl0II
)
,
.CORETSE_AHBo0II
(
CORETSE_AHBo0II
)
)
;
endmodule
