// REVISION    : $Revision: 1.1 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_cnvtxi
(
CORETSE_AHBiO10
,
CORETSE_AHBoi0
,
CORETSE_AHBo11
,
CORETSE_AHBII
,
CORETSE_AHBoI
,
CORETSE_AHBOl
,
CORETSE_AHBIoo0
,
CORETSE_AHBloo0
,
CORETSE_AHBooo0
,
CORETSE_AHBioo0
,
CORETSE_AHBOio0
,
CORETSE_AHBIio0
)
;
input
CORETSE_AHBiO10
;
input
CORETSE_AHBoi0
;
input
[
1
:
0
]
CORETSE_AHBo11
;
input
[
7
:
0
]
CORETSE_AHBII
;
input
CORETSE_AHBoI
;
input
CORETSE_AHBOl
;
input
[
2
:
0
]
CORETSE_AHBIoo0
;
output
[
7
:
0
]
CORETSE_AHBloo0
;
output
CORETSE_AHBooo0
;
output
CORETSE_AHBioo0
;
output
CORETSE_AHBOio0
;
output
[
2
:
0
]
CORETSE_AHBIio0
;
`define CORETSE_AHBIoII  \
# \
1
reg
[
7
:
0
]
CORETSE_AHBlio0
;
reg
[
3
:
0
]
CORETSE_AHBoio0
;
reg
[
3
:
0
]
CORETSE_AHBiio0
;
reg
[
2
:
0
]
CORETSE_AHBOOi0
;
reg
[
1
:
0
]
CORETSE_AHBIOi0
;
reg
[
3
:
0
]
CORETSE_AHBlOi0
;
wire
[
9
:
0
]
CORETSE_AHBoOi0
;
wire
[
2
:
0
]
CORETSE_AHBiOi0
;
reg
[
9
:
0
]
CORETSE_AHBOIi0
;
reg
[
9
:
0
]
CORETSE_AHBIIi0
;
reg
[
9
:
0
]
CORETSE_AHBlIi0
;
reg
[
9
:
0
]
CORETSE_AHBoIi0
;
reg
[
9
:
0
]
CORETSE_AHBiIi0
;
reg
[
9
:
0
]
CORETSE_AHBOli0
;
reg
[
9
:
0
]
CORETSE_AHBIli0
;
reg
[
9
:
0
]
CORETSE_AHBlli0
;
wire
[
9
:
0
]
CORETSE_AHBo0o0
;
reg
[
2
:
0
]
CORETSE_AHBIio0
;
wire
CORETSE_AHBoli0
;
wire
CORETSE_AHBili0
;
reg
CORETSE_AHBOio0
;
reg
[
2
:
0
]
CORETSE_AHBO0i0
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBlio0
<=
`CORETSE_AHBIoII
8
'h
00
;
else
CORETSE_AHBlio0
<=
`CORETSE_AHBIoII
CORETSE_AHBII
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBoio0
<=
`CORETSE_AHBIoII
4
'h
0
;
else
CORETSE_AHBoio0
<=
`CORETSE_AHBIoII
CORETSE_AHBlio0
[
3
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBiio0
<=
`CORETSE_AHBIoII
4
'h
0
;
else
CORETSE_AHBiio0
<=
`CORETSE_AHBIoII
CORETSE_AHBoio0
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBOOi0
<=
`CORETSE_AHBIoII
3
'h
0
;
else
CORETSE_AHBOOi0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBOOi0
[
1
:
0
]
,
CORETSE_AHBoI
}
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBIOi0
<=
`CORETSE_AHBIoII
2
'h
0
;
else
CORETSE_AHBIOi0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBIOi0
[
0
]
,
CORETSE_AHBOl
}
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBlOi0
<=
`CORETSE_AHBIoII
4
'h
0
;
else
if
(
~
(
~
CORETSE_AHBOOi0
[
1
]
&
CORETSE_AHBOOi0
[
0
]
&
CORETSE_AHBlOi0
[
0
]
&
(
CORETSE_AHBo11
!=
2
'b
10
)
)
)
CORETSE_AHBlOi0
<=
`CORETSE_AHBIoII
CORETSE_AHBlOi0
+
4
'h
1
;
end
assign
CORETSE_AHBoOi0
=
(
{
10
{
CORETSE_AHBo11
==
2
'b
10
}
}
&
{
CORETSE_AHBIOi0
[
0
]
,
CORETSE_AHBOOi0
[
0
]
,
CORETSE_AHBlio0
}
)
|
(
{
10
{
(
CORETSE_AHBo11
!=
2
'b
10
)
&
CORETSE_AHBlOi0
[
0
]
}
}
&
{
(
CORETSE_AHBIOi0
[
1
]
|
CORETSE_AHBIOi0
[
0
]
)
,
(
CORETSE_AHBOOi0
[
1
]
|
CORETSE_AHBOOi0
[
0
]
)
,
CORETSE_AHBlio0
[
3
:
0
]
,
CORETSE_AHBoio0
[
3
:
0
]
}
)
;
assign
CORETSE_AHBiOi0
=
(
{
3
{
(
CORETSE_AHBo11
==
2
'b
10
)
}
}
&
CORETSE_AHBlOi0
[
2
:
0
]
)
|
(
{
3
{
(
CORETSE_AHBo11
!=
2
'b
10
)
}
}
&
CORETSE_AHBlOi0
[
3
:
1
]
)
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
begin
CORETSE_AHBOIi0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBIIi0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBlIi0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBoIi0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBiIi0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBOli0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBIli0
<=
`CORETSE_AHBIoII
10
'h
000
;
CORETSE_AHBlli0
<=
`CORETSE_AHBIoII
10
'h
000
;
end
else
case
(
CORETSE_AHBiOi0
)
3
'h
0
:
CORETSE_AHBOIi0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
1
:
CORETSE_AHBIIi0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
2
:
CORETSE_AHBlIi0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
3
:
CORETSE_AHBoIi0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
4
:
CORETSE_AHBiIi0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
5
:
CORETSE_AHBOli0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
6
:
CORETSE_AHBIli0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
3
'h
7
:
CORETSE_AHBlli0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
default
:
CORETSE_AHBOIi0
<=
`CORETSE_AHBIoII
CORETSE_AHBoOi0
;
endcase
end
assign
CORETSE_AHBoli0
=
(
(
(
CORETSE_AHBo11
==
2
'b
10
)
&
(
CORETSE_AHBOOi0
[
0
]
==
1
'b
1
)
)
|
(
(
CORETSE_AHBo11
!=
2
'b
10
)
&
(
CORETSE_AHBOOi0
[
1
]
==
1
'b
1
)
)
|
(
~
CORETSE_AHBOio0
&
~
(
|
CORETSE_AHBO0i0
)
&
CORETSE_AHBlOi0
[
0
]
)
&
~
(
|
CORETSE_AHBOOi0
)
)
;
assign
CORETSE_AHBili0
=
(
(
(
CORETSE_AHBo11
==
2
'b
10
)
&
(
CORETSE_AHBOOi0
[
1
:
0
]
==
2
'b
10
)
)
|
(
(
CORETSE_AHBo11
!=
2
'b
10
)
&
(
CORETSE_AHBOOi0
[
2
:
1
]
==
2
'b
10
)
)
|
(
CORETSE_AHBOio0
&
CORETSE_AHBO0i0
[
0
]
)
)
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBOio0
<=
`CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBoli0
)
CORETSE_AHBOio0
<=
`CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBili0
)
CORETSE_AHBOio0
<=
`CORETSE_AHBIoII
1
'b
0
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBO0i0
<=
`CORETSE_AHBIoII
3
'h
0
;
else
CORETSE_AHBO0i0
<=
`CORETSE_AHBIoII
{
CORETSE_AHBO0i0
[
1
:
0
]
,
CORETSE_AHBOio0
}
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBiO10
)
begin
if
(
CORETSE_AHBiO10
)
CORETSE_AHBIio0
<=
`CORETSE_AHBIoII
3
'h
0
;
else
if
(
~
CORETSE_AHBOio0
&
CORETSE_AHBoli0
&
(
CORETSE_AHBo11
==
2
'b
10
)
)
CORETSE_AHBIio0
<=
`CORETSE_AHBIoII
CORETSE_AHBiOi0
;
else
if
(
~
CORETSE_AHBOio0
&
CORETSE_AHBoli0
&
(
CORETSE_AHBo11
!=
2
'b
10
)
)
CORETSE_AHBIio0
<=
`CORETSE_AHBIoII
CORETSE_AHBiOi0
+
3
'h
5
;
end
assign
CORETSE_AHBo0o0
=
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
0
)
}
}
&
CORETSE_AHBOIi0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
1
)
}
}
&
CORETSE_AHBIIi0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
2
)
}
}
&
CORETSE_AHBlIi0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
3
)
}
}
&
CORETSE_AHBoIi0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
4
)
}
}
&
CORETSE_AHBiIi0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
5
)
}
}
&
CORETSE_AHBOli0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
6
)
}
}
&
CORETSE_AHBIli0
|
{
10
{
(
CORETSE_AHBIoo0
==
3
'h
7
)
}
}
&
CORETSE_AHBlli0
;
assign
CORETSE_AHBloo0
=
CORETSE_AHBo0o0
[
7
:
0
]
;
assign
CORETSE_AHBooo0
=
CORETSE_AHBo0o0
[
8
]
;
assign
CORETSE_AHBioo0
=
CORETSE_AHBo0o0
[
9
]
;
endmodule
