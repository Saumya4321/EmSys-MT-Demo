// REVISION    : $Revision: 1.7 $
//         Mentor Graphics Corporation Proprietary and Confidential
//         Copyright Mentor Graphics Corporation and Licensors 2004
`include "include.v"
module
dmatx
#
(
parameter
CORETSE_AHBoOI
=
0
)
(
CORETSE_AHBI01l
,
HREADY
,
HRESP
,
HRDATA
,
CORETSE_AHBl1Il
,
HCLK
,
CORETSE_AHBl01l
,
HTRANS
,
HADDR
,
HWRITE
,
HWDATA
,
CORETSE_AHBi00l
,
CORETSE_AHBOo0l
,
CORETSE_AHBo10l
,
CORETSE_AHBil0l
,
CORETSE_AHBioll
,
CORETSE_AHBOill
,
CORETSE_AHBol1l
,
CORETSE_AHBI10l
,
CORETSE_AHBII0l
,
CORETSE_AHBiIll
,
CORETSE_AHBOlll
,
CORETSE_AHBIlll
,
CORETSE_AHBllll
,
CORETSE_AHBolll
,
CORETSE_AHBO0ll
,
CORETSE_AHBI0ll
,
CORETSE_AHBl0ll
,
CORETSE_AHBo0ll
,
CORETSE_AHBi0ll
,
CORETSE_AHBO1ll
)
;
input
CORETSE_AHBI01l
;
input
HREADY
;
input
[
1
:
0
]
HRESP
;
input
[
31
:
0
]
HRDATA
;
input
CORETSE_AHBl1Il
;
input
HCLK
;
output
CORETSE_AHBl01l
;
output
[
1
:
0
]
HTRANS
;
output
[
31
:
2
]
HADDR
;
output
HWRITE
;
output
[
31
:
0
]
HWDATA
;
input
[
31
:
2
]
CORETSE_AHBI10l
;
output
CORETSE_AHBi00l
;
output
CORETSE_AHBOo0l
;
output
[
31
:
2
]
CORETSE_AHBo10l
;
input
CORETSE_AHBioll
;
input
CORETSE_AHBOill
;
input
CORETSE_AHBol1l
;
output
CORETSE_AHBII0l
;
output
[
7
:
0
]
CORETSE_AHBil0l
;
output
CORETSE_AHBiIll
;
output
CORETSE_AHBOlll
;
output
CORETSE_AHBIlll
;
output
[
31
:
0
]
CORETSE_AHBllll
;
output
[
1
:
0
]
CORETSE_AHBolll
;
output
CORETSE_AHBO0ll
;
output
CORETSE_AHBI0ll
;
output
[
1
:
0
]
CORETSE_AHBl0ll
;
output
CORETSE_AHBo0ll
;
input
CORETSE_AHBi0ll
;
input
CORETSE_AHBO1ll
;
`define CORETSE_AHBi01l  \
2 \
'b \
00
`define CORETSE_AHBO11l  \
2 \
'b \
01
`define CORETSE_AHBI11l  \
2 \
'b \
11
`define CORETSE_AHBl11l  \
2 \
'b \
10
`define CORETSE_AHBo11l  \
1 \
'b \
0
`define CORETSE_AHBi11l  \
1 \
'b \
1
`define CORETSE_AHBOo1l  \
{ \
1 \
'b \
0 \
, \
`CORETSE_AHBIo1l \
}
`define CORETSE_AHBlo1l  \
{ \
1 \
'b \
1 \
, \
`CORETSE_AHBIo1l \
}
`define CORETSE_AHBoo1l  \
{ \
1 \
'b \
1 \
, \
`CORETSE_AHBio1l \
}
`define CORETSE_AHBOi1l  \
{ \
1 \
'b \
1 \
, \
`CORETSE_AHBIi1l \
}
`define CORETSE_AHBli1l  \
{ \
1 \
'b \
1 \
, \
`CORETSE_AHBoi1l \
}
reg
[
1
:
0
]
CORETSE_AHBOOol
,
CORETSE_AHBIOol
;
reg
CORETSE_AHBII0l
;
reg
[
7
:
0
]
CORETSE_AHBil0l
,
CORETSE_AHBIiol
;
reg
CORETSE_AHBliol
;
reg
CORETSE_AHBOo0l
;
reg
[
31
:
2
]
CORETSE_AHBo10l
;
reg
[
1
:
0
]
CORETSE_AHBiOol
;
reg
[
31
:
2
]
CORETSE_AHBOIol
;
reg
CORETSE_AHBIIol
;
reg
[
15
:
0
]
CORETSE_AHBoiol
;
reg
[
4
:
0
]
CORETSE_AHBiiol
;
reg
[
31
:
2
]
CORETSE_AHBlIol
;
reg
[
31
:
2
]
CORETSE_AHBiIol
;
reg
[
15
:
0
]
CORETSE_AHBOlol
;
reg
[
15
:
0
]
CORETSE_AHBIlol
;
reg
CORETSE_AHBllol
;
reg
CORETSE_AHBolol
;
reg
CORETSE_AHBilol
;
reg
[
31
:
0
]
CORETSE_AHBO0ol
;
reg
[
2
:
0
]
CORETSE_AHBI0ol
,
CORETSE_AHBl0ol
;
reg
CORETSE_AHBo0ol
;
reg
CORETSE_AHBi0ol
;
wire
CORETSE_AHBO1ol
;
reg
HWRITE
;
reg
[
31
:
0
]
HWDATA
;
reg
[
31
:
2
]
HADDR
,
CORETSE_AHBI1ol
;
reg
[
15
:
0
]
CORETSE_AHBl1ol
,
CORETSE_AHBo1ol
;
reg
CORETSE_AHBOOil
;
reg
CORETSE_AHBIOil
;
reg
CORETSE_AHBOlll
;
reg
CORETSE_AHBIlll
;
reg
CORETSE_AHBiIll
;
reg
[
1
:
0
]
CORETSE_AHBolll
;
reg
[
31
:
0
]
CORETSE_AHBllll
;
wire
CORETSE_AHBlOil
;
assign
CORETSE_AHBi00l
=
CORETSE_AHBO1ol
;
assign
CORETSE_AHBlOil
=
CORETSE_AHBII0l
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBoOil
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBII0l
<=
0
;
CORETSE_AHBil0l
<=
0
;
end
else
begin
CORETSE_AHBII0l
<=
(
CORETSE_AHBII0l
||
CORETSE_AHBioll
)
&&
CORETSE_AHBliol
&&
!
CORETSE_AHBOill
;
CORETSE_AHBil0l
<=
CORETSE_AHBIiol
-
{
7
'h
00
,
(
CORETSE_AHBol1l
&&
|
CORETSE_AHBil0l
)
}
;
end
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBOool
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBOOol
<=
`CORETSE_AHBi01l
;
CORETSE_AHBlIol
<=
0
;
CORETSE_AHBoiol
<=
0
;
CORETSE_AHBIIol
<=
0
;
CORETSE_AHBiiol
<=
0
;
CORETSE_AHBOIol
<=
0
;
CORETSE_AHBiOol
<=
0
;
end
else
begin
CORETSE_AHBOOol
<=
CORETSE_AHBIOol
;
if
(
HREADY
)
if
(
CORETSE_AHBOOol
==
`CORETSE_AHBO11l
)
CORETSE_AHBiOol
<=
CORETSE_AHBl1ol
+
1
;
else
CORETSE_AHBiOol
<=
0
;
case
(
CORETSE_AHBiOol
)
2
'b
11
:
CORETSE_AHBlIol
<=
HRDATA
[
31
:
2
]
;
2
'b
10
:
begin
CORETSE_AHBoiol
<=
HRDATA
[
15
:
0
]
;
CORETSE_AHBiiol
<=
HRDATA
[
20
:
16
]
;
CORETSE_AHBIIol
<=
HRDATA
[
31
]
;
end
2
'b
01
:
CORETSE_AHBOIol
<=
HRDATA
[
31
:
2
]
;
endcase
end
end
always
@
(
*
)
begin
:
CORETSE_AHBIool
CORETSE_AHBIOol
=
CORETSE_AHBOOol
;
CORETSE_AHBliol
=
1
;
CORETSE_AHBOo0l
=
0
;
CORETSE_AHBIiol
=
CORETSE_AHBil0l
;
CORETSE_AHBo10l
=
CORETSE_AHBI10l
;
if
(
CORETSE_AHBO1ol
)
begin
CORETSE_AHBIOol
=
`CORETSE_AHBi01l
;
CORETSE_AHBliol
=
0
;
end
else
case
(
CORETSE_AHBOOol
)
`CORETSE_AHBi01l
:
begin
if
(
CORETSE_AHBlOil
)
CORETSE_AHBIOol
=
`CORETSE_AHBO11l
;
else
CORETSE_AHBIOol
=
`CORETSE_AHBi01l
;
end
`CORETSE_AHBO11l
:
begin
if
(
CORETSE_AHBi0ol
)
if
(
(
CORETSE_AHBiOol
==
2
'b
10
)
?
HRDATA
[
31
]
:
CORETSE_AHBIIol
)
begin
CORETSE_AHBliol
=
0
;
CORETSE_AHBOo0l
=
1
;
CORETSE_AHBIOol
=
`CORETSE_AHBi01l
;
end
else
CORETSE_AHBIOol
=
`CORETSE_AHBI11l
;
end
`CORETSE_AHBI11l
:
begin
if
(
CORETSE_AHBi0ol
)
CORETSE_AHBIOol
=
`CORETSE_AHBl11l
;
end
`CORETSE_AHBl11l
:
begin
if
(
CORETSE_AHBi0ol
)
begin
CORETSE_AHBIiol
=
CORETSE_AHBil0l
+
1
;
if
(
CORETSE_AHBlOil
)
begin
CORETSE_AHBIOol
=
`CORETSE_AHBO11l
;
end
else
begin
CORETSE_AHBIOol
=
`CORETSE_AHBi01l
;
end
end
end
endcase
if
(
CORETSE_AHBI01l
&&
HREADY
&&
CORETSE_AHBIOol
==
`CORETSE_AHBl11l
)
CORETSE_AHBo10l
=
CORETSE_AHBOIol
;
end
always
@
(
CORETSE_AHBIOol
or
CORETSE_AHBOOol
or
CORETSE_AHBiOol
or
CORETSE_AHBO1ll
or
CORETSE_AHBI10l
or
CORETSE_AHBl1ol
or
CORETSE_AHBoiol
or
CORETSE_AHBlIol
or
HRDATA
or
CORETSE_AHBi0ll
)
begin
:
CORETSE_AHBlool
case
(
CORETSE_AHBIOol
)
`CORETSE_AHBO11l
:
begin
CORETSE_AHBIlol
=
16
'h
0002
;
CORETSE_AHBilol
=
0
;
CORETSE_AHBllol
=
1
;
CORETSE_AHBiIol
=
CORETSE_AHBI10l
;
end
`CORETSE_AHBI11l
:
begin
CORETSE_AHBilol
=
0
;
CORETSE_AHBIlol
=
(
CORETSE_AHBiOol
==
2
'b
10
)
?
HRDATA
[
15
:
0
]
-
1
:
CORETSE_AHBoiol
-
1
;
CORETSE_AHBllol
=
!
CORETSE_AHBO1ll
&&
CORETSE_AHBi0ll
;
CORETSE_AHBiIol
=
CORETSE_AHBlIol
;
end
`CORETSE_AHBl11l
:
begin
CORETSE_AHBIlol
=
CORETSE_AHBl1ol
+
16
'h
0004
;
CORETSE_AHBilol
=
1
;
CORETSE_AHBllol
=
1
;
CORETSE_AHBiIol
=
CORETSE_AHBI10l
+
1
;
end
default
:
begin
CORETSE_AHBIlol
=
0
;
CORETSE_AHBilol
=
0
;
CORETSE_AHBllol
=
0
;
CORETSE_AHBiIol
=
0
;
end
endcase
case
(
CORETSE_AHBOOol
)
`CORETSE_AHBO11l
:
begin
CORETSE_AHBOlol
=
16
'h
FFFF
;
CORETSE_AHBolol
=
~|
CORETSE_AHBl1ol
;
CORETSE_AHBO0ol
=
0
;
end
`CORETSE_AHBI11l
:
begin
CORETSE_AHBOlol
=
16
'h
FFFC
;
CORETSE_AHBolol
=
~|
CORETSE_AHBl1ol
[
15
:
2
]
||
!
CORETSE_AHBi0ll
;
CORETSE_AHBO0ol
=
HRDATA
;
end
`CORETSE_AHBl11l
:
begin
CORETSE_AHBOlol
=
0
;
CORETSE_AHBolol
=
1
;
CORETSE_AHBO0ol
[
31
]
=
1
;
CORETSE_AHBO0ol
[
30
:
0
]
=
0
;
end
default
:
begin
CORETSE_AHBOlol
=
0
;
CORETSE_AHBolol
=
1
;
CORETSE_AHBO0ol
=
0
;
end
endcase
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBoool
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBI0ol
<=
`CORETSE_AHBOo1l
;
CORETSE_AHBo0ol
<=
0
;
HADDR
<=
0
;
HWRITE
<=
0
;
HWDATA
<=
0
;
CORETSE_AHBl1ol
<=
0
;
end
else
begin
CORETSE_AHBI0ol
<=
CORETSE_AHBl0ol
;
CORETSE_AHBo0ol
<=
HREADY
?
CORETSE_AHBI0ol
[
1
]
:
CORETSE_AHBo0ol
;
HWDATA
<=
HREADY
?
CORETSE_AHBO0ol
:
HWDATA
;
HWRITE
<=
HREADY
?
CORETSE_AHBilol
:
HWRITE
;
HADDR
<=
CORETSE_AHBI1ol
;
CORETSE_AHBl1ol
<=
CORETSE_AHBo1ol
;
end
end
assign
CORETSE_AHBO1ol
=
CORETSE_AHBo0ol
&&
HREADY
&&
(
HRESP
!=
`CORETSE_AHBiool
)
;
always
@
(
HREADY
or
CORETSE_AHBI0ol
or
CORETSE_AHBI01l
or
HADDR
or
CORETSE_AHBllol
or
CORETSE_AHBolol
or
CORETSE_AHBiIol
or
CORETSE_AHBIlol
or
CORETSE_AHBOlol
or
CORETSE_AHBl1ol
)
begin
:
CORETSE_AHBOiol
CORETSE_AHBl0ol
=
CORETSE_AHBI0ol
;
CORETSE_AHBI1ol
=
HADDR
;
CORETSE_AHBo1ol
=
CORETSE_AHBl1ol
;
CORETSE_AHBi0ol
=
0
;
if
(
HREADY
)
case
(
CORETSE_AHBI0ol
)
`CORETSE_AHBOo1l
:
if
(
CORETSE_AHBllol
)
begin
CORETSE_AHBl0ol
=
CORETSE_AHBI01l
?
`CORETSE_AHBOi1l
:
`CORETSE_AHBlo1l
;
CORETSE_AHBI1ol
=
CORETSE_AHBiIol
;
CORETSE_AHBo1ol
=
CORETSE_AHBIlol
;
end
`CORETSE_AHBlo1l
:
CORETSE_AHBl0ol
=
CORETSE_AHBI01l
?
`CORETSE_AHBOi1l
:
`CORETSE_AHBlo1l
;
`CORETSE_AHBOi1l
,
`CORETSE_AHBli1l
:
begin
CORETSE_AHBI1ol
=
HADDR
+
1
;
CORETSE_AHBo1ol
=
CORETSE_AHBl1ol
+
CORETSE_AHBOlol
;
if
(
CORETSE_AHBolol
)
begin
CORETSE_AHBi0ol
=
1
;
if
(
CORETSE_AHBllol
&&
CORETSE_AHBI01l
)
begin
CORETSE_AHBI1ol
=
CORETSE_AHBiIol
;
CORETSE_AHBo1ol
=
CORETSE_AHBIlol
;
CORETSE_AHBl0ol
=
`CORETSE_AHBOi1l
;
end
else
CORETSE_AHBl0ol
=
`CORETSE_AHBOo1l
;
end
else
if
(
!
CORETSE_AHBI01l
)
CORETSE_AHBl0ol
=
`CORETSE_AHBlo1l
;
else
if
(
~|
CORETSE_AHBI1ol
[
9
:
2
]
)
CORETSE_AHBl0ol
=
`CORETSE_AHBOi1l
;
else
CORETSE_AHBl0ol
=
`CORETSE_AHBli1l
;
end
default
:
begin
CORETSE_AHBl0ol
=
`CORETSE_AHBOo1l
;
end
endcase
end
assign
HTRANS
=
CORETSE_AHBI0ol
[
1
:
0
]
;
assign
CORETSE_AHBl01l
=
CORETSE_AHBI0ol
[
2
]
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBiOil
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBOOil
<=
0
;
CORETSE_AHBIOil
<=
0
;
CORETSE_AHBiIll
<=
0
;
CORETSE_AHBOlll
<=
0
;
CORETSE_AHBIlll
<=
0
;
CORETSE_AHBolll
<=
0
;
CORETSE_AHBllll
<=
0
;
end
else
begin
if
(
HREADY
&&
CORETSE_AHBI0ol
[
1
]
)
begin
CORETSE_AHBOOil
<=
(
CORETSE_AHBOOol
==
`CORETSE_AHBI11l
)
;
CORETSE_AHBIOil
<=
(
CORETSE_AHBOOol
==
`CORETSE_AHBI11l
)
&&
!
CORETSE_AHBOOil
;
end
if
(
CORETSE_AHBOOil
&&
CORETSE_AHBo0ol
&&
HREADY
)
begin
CORETSE_AHBiIll
<=
1
;
CORETSE_AHBOlll
<=
CORETSE_AHBIOil
;
CORETSE_AHBIlll
<=
CORETSE_AHBOOil
&&
(
CORETSE_AHBOOol
!=
`CORETSE_AHBI11l
)
;
CORETSE_AHBolll
<=
CORETSE_AHBOOil
&&
(
CORETSE_AHBOOol
!=
`CORETSE_AHBI11l
)
?
~
CORETSE_AHBl1ol
[
1
:
0
]
:
0
;
CORETSE_AHBllll
<=
HRDATA
;
end
else
begin
CORETSE_AHBiIll
<=
0
;
CORETSE_AHBOlll
<=
0
;
CORETSE_AHBIlll
<=
0
;
CORETSE_AHBolll
<=
0
;
CORETSE_AHBllll
<=
0
;
end
end
end
assign
CORETSE_AHBO0ll
=
CORETSE_AHBiiol
[
0
]
;
assign
CORETSE_AHBI0ll
=
CORETSE_AHBiiol
[
1
]
;
assign
CORETSE_AHBl0ll
=
CORETSE_AHBiiol
[
3
:
2
]
;
assign
CORETSE_AHBo0ll
=
CORETSE_AHBiiol
[
4
]
;
endmodule
