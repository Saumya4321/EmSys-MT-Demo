// REVISION    : $Revision: 1.1 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
r10b8b
(
CORETSE_AHBIoIOI
,
CORETSE_AHBOloi
,
CORETSE_AHBOo1
,
CORETSE_AHBo0o
,
CORETSE_AHBo0oi
,
CORETSE_AHBO0oi
,
CORETSE_AHBi0oi
)
;
input
[
9
:
0
]
CORETSE_AHBIoIOI
;
input
CORETSE_AHBOloi
;
input
CORETSE_AHBOo1
;
output
[
7
:
0
]
CORETSE_AHBo0o
;
output
[
2
:
0
]
CORETSE_AHBo0oi
;
output
CORETSE_AHBO0oi
;
output
CORETSE_AHBi0oi
;
parameter
CORETSE_AHBIoII
=
1
;
wire
[
9
:
0
]
CORETSE_AHBlii1I
;
wire
[
5
:
0
]
CORETSE_AHBoii1I
;
wire
[
3
:
0
]
CORETSE_AHBiii1I
;
reg
[
4
:
0
]
CORETSE_AHBOOOoI
;
reg
CORETSE_AHBIOOoI
;
reg
[
1
:
0
]
CORETSE_AHBlOOoI
;
reg
CORETSE_AHBoOOoI
;
reg
[
1
:
0
]
CORETSE_AHBiOOoI
;
reg
[
2
:
0
]
CORETSE_AHBOIOoI
;
reg
CORETSE_AHBIIOoI
,
CORETSE_AHBlIOoI
;
reg
[
1
:
0
]
CORETSE_AHBoIOoI
;
reg
[
2
:
0
]
CORETSE_AHBiIOoI
;
wire
[
7
:
0
]
CORETSE_AHBOlOoI
;
wire
CORETSE_AHBIlOoI
;
reg
[
2
:
0
]
CORETSE_AHBllOoI
;
reg
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
;
wire
CORETSE_AHBO0OoI
;
reg
CORETSE_AHBI0OoI
;
reg
[
2
:
0
]
CORETSE_AHBl0OoI
;
reg
[
7
:
0
]
CORETSE_AHBo0OoI
;
assign
CORETSE_AHBlii1I
=
{
CORETSE_AHBIoIOI
[
6
]
,
CORETSE_AHBIoIOI
[
7
]
,
CORETSE_AHBIoIOI
[
8
]
,
CORETSE_AHBIoIOI
[
9
]
,
CORETSE_AHBIoIOI
[
0
]
,
CORETSE_AHBIoIOI
[
1
]
,
CORETSE_AHBIoIOI
[
2
]
,
CORETSE_AHBIoIOI
[
3
]
,
CORETSE_AHBIoIOI
[
4
]
,
CORETSE_AHBIoIOI
[
5
]
}
;
assign
CORETSE_AHBoii1I
=
CORETSE_AHBlii1I
[
5
:
0
]
;
always
@
(
CORETSE_AHBlii1I
[
5
:
0
]
)
case
(
{
CORETSE_AHBlii1I
[
5
]
,
CORETSE_AHBlii1I
[
4
]
,
CORETSE_AHBlii1I
[
3
]
,
CORETSE_AHBlii1I
[
2
]
,
CORETSE_AHBlii1I
[
1
]
,
CORETSE_AHBlii1I
[
0
]
}
)
6
'b
100111
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00000_1_10_0_00
;
6
'b
011000
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00000_1_11_0_00
;
6
'b
011101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00001_1_10_0_00
;
6
'b
100010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00001_1_11_0_00
;
6
'b
101101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00010_1_10_0_00
;
6
'b
010010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00010_1_11_0_00
;
6
'b
110001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00011_1_00_1_00
;
6
'b
110101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00100_1_10_0_00
;
6
'b
001010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00100_1_11_0_00
;
6
'b
101001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00101_1_00_1_00
;
6
'b
011001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00110_1_00_1_00
;
6
'b
111000
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00111_1_10_1_00
;
6
'b
000111
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00111_1_11_1_00
;
6
'b
111001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01000_1_10_0_00
;
6
'b
000110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01000_1_11_0_00
;
6
'b
100101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01001_1_00_1_00
;
6
'b
010101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01010_1_00_1_00
;
6
'b
110100
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01011_1_00_1_01
;
6
'b
001101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01100_1_00_1_00
;
6
'b
101100
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01101_1_00_1_01
;
6
'b
011100
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01110_1_00_1_01
;
6
'b
010111
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01111_1_10_0_00
;
6
'b
101000
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
01111_1_11_0_00
;
6
'b
011011
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10000_1_10_0_00
;
6
'b
100100
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10000_1_11_0_00
;
6
'b
100011
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10001_1_00_1_10
;
6
'b
010011
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10010_1_00_1_10
;
6
'b
110010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10011_1_00_1_00
;
6
'b
001011
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10100_1_00_1_10
;
6
'b
101010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10101_1_00_1_00
;
6
'b
011010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10110_1_00_1_00
;
6
'b
111010
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10111_1_10_0_00
;
6
'b
000101
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
10111_1_11_0_00
;
6
'b
110011
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11000_1_10_0_00
;
6
'b
001100
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11000_1_11_0_00
;
6
'b
100110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11001_1_00_1_00
;
6
'b
010110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11010_1_00_1_00
;
6
'b
110110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11011_1_10_0_00
;
6
'b
001001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11011_1_11_0_00
;
6
'b
001110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11100_1_00_1_00
;
6
'b
101110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11101_1_10_0_00
;
6
'b
010001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11101_1_11_0_00
;
6
'b
011110
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11110_1_10_0_00
;
6
'b
100001
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11110_1_11_0_00
;
6
'b
101011
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11111_1_10_0_00
;
6
'b
010100
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
11111_1_11_0_00
;
default
:
{
CORETSE_AHBOOOoI
,
CORETSE_AHBIOOoI
,
CORETSE_AHBlOOoI
,
CORETSE_AHBoOOoI
,
CORETSE_AHBiOOoI
}
=
11
'b
00000_0_00_0_00
;
endcase
assign
CORETSE_AHBiii1I
=
CORETSE_AHBlii1I
[
9
:
6
]
;
always
@
(
CORETSE_AHBlii1I
[
9
:
6
]
)
case
(
{
CORETSE_AHBlii1I
[
9
]
,
CORETSE_AHBlii1I
[
8
]
,
CORETSE_AHBlii1I
[
7
]
,
CORETSE_AHBlii1I
[
6
]
}
)
4
'b
1011
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
000_1_11__000_0
;
4
'b
0100
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
000_1_10__000_0
;
4
'b
1001
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
001_1_00__000_1
;
4
'b
0101
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
010_1_00__000_1
;
4
'b
0011
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
011_1_10__000_1
;
4
'b
1100
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
011_1_11__000_1
;
4
'b
0010
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
100_1_10__000_0
;
4
'b
1101
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
100_1_11__000_0
;
4
'b
1010
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
101_1_00__000_1
;
4
'b
0110
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
110_1_00__000_1
;
4
'b
0001
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
111_1_10__100_0
;
4
'b
1110
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
111_1_11__100_0
;
4
'b
0111
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
111_1_00__110_0
;
4
'b
1000
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
111_1_00__101_0
;
default
:
{
CORETSE_AHBOIOoI
,
CORETSE_AHBIIOoI
,
CORETSE_AHBoIOoI
,
CORETSE_AHBiIOoI
,
CORETSE_AHBlIOoI
}
=
10
'b
000_0_00__000_0
;
endcase
assign
CORETSE_AHBOlOoI
=
{
CORETSE_AHBOIOoI
,
CORETSE_AHBOOOoI
}
;
assign
CORETSE_AHBIlOoI
=
CORETSE_AHBIOOoI
&
CORETSE_AHBIIOoI
&
(
(
CORETSE_AHBOloi
&
CORETSE_AHBlOOoI
[
1
]
)
==
CORETSE_AHBlOOoI
[
0
]
)
&
(
CORETSE_AHBiIOoI
[
1
]
|
CORETSE_AHBiIOoI
[
0
]
|
(
(
CORETSE_AHBoIOoI
[
1
]
&
(
CORETSE_AHBOloi
^
CORETSE_AHBoOOoI
)
)
==
CORETSE_AHBoIOoI
[
0
]
)
)
&
(
~
CORETSE_AHBiIOoI
[
1
]
&
(
~
CORETSE_AHBiOOoI
[
1
]
|
CORETSE_AHBOloi
|
~
CORETSE_AHBiIOoI
[
2
]
)
|
CORETSE_AHBiIOoI
[
1
]
&
CORETSE_AHBiOOoI
[
1
]
&
~
CORETSE_AHBOloi
&
CORETSE_AHBiIOoI
[
2
]
)
&
(
~
CORETSE_AHBiIOoI
[
0
]
&
(
~
CORETSE_AHBiOOoI
[
0
]
|
~
CORETSE_AHBOloi
|
~
CORETSE_AHBiIOoI
[
2
]
)
|
CORETSE_AHBiIOoI
[
0
]
&
CORETSE_AHBiOOoI
[
0
]
&
CORETSE_AHBOloi
&
CORETSE_AHBiIOoI
[
2
]
)
;
assign
CORETSE_AHBi0oi
=
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
11_0111_1100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
00_0111_1100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_1111_1100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0011_1100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0101_1100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0110_1100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0111_0100
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0111_1000
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0111_1110
)
|
~
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
01_0111_1101
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
00_1000_0011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
11_1000_0011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_0000_0011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1100_0011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1010_0011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1001_0011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1000_1011
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1000_0111
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1000_0001
)
|
CORETSE_AHBOloi
&
(
CORETSE_AHBIoIOI
==
10
'b
10_1000_0010
)
;
always
@
(
CORETSE_AHBlii1I
)
casex
(
{
CORETSE_AHBlii1I
[
9
]
,
CORETSE_AHBlii1I
[
8
]
,
CORETSE_AHBlii1I
[
7
]
,
CORETSE_AHBlii1I
[
6
]
,
CORETSE_AHBlii1I
[
5
]
,
CORETSE_AHBlii1I
[
4
]
,
CORETSE_AHBlii1I
[
3
]
,
CORETSE_AHBlii1I
[
2
]
,
CORETSE_AHBlii1I
[
1
]
,
CORETSE_AHBlii1I
[
0
]
}
)
10
'b
10_0011_0110
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
000_1_0
;
10
'b
01_1100_1001
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
000_1_1
;
10
'b
10_0010_1110
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
010_1_0
;
10
'b
01_1101_0001
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
010_1_1
;
10
'b
10_0011_1010
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
011_1_0
;
10
'b
01_1100_0101
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
011_1_1
;
10
'b
10_1000_1111
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
100_1_0
;
10
'b
01_0111_0000
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
100_1_1
;
10
'b
10_0100_1111
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
100_1_0
;
10
'b
01_1011_0000
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
100_1_1
;
10
'b
10_0001_1110
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
111_1_0
;
10
'b
01_1110_0001
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
111_1_1
;
default
:
{
CORETSE_AHBllOoI
,
CORETSE_AHBolOoI
,
CORETSE_AHBilOoI
}
=
5
'b
001_0_0
;
endcase
assign
CORETSE_AHBO0OoI
=
~
CORETSE_AHBOo1
&
CORETSE_AHBolOoI
|
CORETSE_AHBOo1
&
CORETSE_AHBolOoI
&
(
CORETSE_AHBilOoI
==
CORETSE_AHBOloi
)
;
always
@
(
CORETSE_AHBO0OoI
or
CORETSE_AHBIlOoI
or
CORETSE_AHBOlOoI
or
CORETSE_AHBllOoI
or
CORETSE_AHBoOOoI
or
CORETSE_AHBlIOoI
)
begin
casex
(
{
CORETSE_AHBO0OoI
,
CORETSE_AHBIlOoI
,
CORETSE_AHBllOoI
}
)
5
'b
0_0_xxx
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
12
'b
001_00000000_0
;
5
'b
0_1_xxx
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
{
3
'b
101
,
CORETSE_AHBOlOoI
,
CORETSE_AHBoOOoI
^
CORETSE_AHBlIOoI
}
;
5
'b
1_0_000
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
{
CORETSE_AHBllOoI
,
8
'h
fb
,
1
'b
0
}
;
5
'b
1_0_010
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
{
CORETSE_AHBllOoI
,
8
'h
fd
,
1
'b
0
}
;
5
'b
1_0_011
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
{
CORETSE_AHBllOoI
,
8
'h
f7
,
1
'b
0
}
;
5
'b
1_0_100
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
{
CORETSE_AHBllOoI
,
8
'h
bc
,
1
'b
1
}
;
5
'b
1_0_111
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
{
CORETSE_AHBllOoI
,
8
'h
fe
,
1
'b
0
}
;
5
'b
1_1_xxx
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
12
'b
001_00000000_0
;
default
:
{
CORETSE_AHBl0OoI
,
CORETSE_AHBo0OoI
,
CORETSE_AHBI0OoI
}
=
12
'b
001_00000000_0
;
endcase
end
assign
CORETSE_AHBo0o
=
CORETSE_AHBo0OoI
;
assign
CORETSE_AHBo0oi
=
CORETSE_AHBl0OoI
;
reg
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
;
always
@
(
CORETSE_AHBlii1I
[
5
:
0
]
)
case
(
{
CORETSE_AHBlii1I
[
5
]
,
CORETSE_AHBlii1I
[
4
]
,
CORETSE_AHBlii1I
[
3
]
,
CORETSE_AHBlii1I
[
2
]
,
CORETSE_AHBlii1I
[
1
]
,
CORETSE_AHBlii1I
[
0
]
}
)
6
'b
000000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
000111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
001000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
001001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
001010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
001011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
001100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
001101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
001110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
001111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
010000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
010001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
010010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
010011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
010100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
010101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
010110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
010111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
011000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
011001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
011010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
011011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
011100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
011101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
011110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
011111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
100000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
100001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
100010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
100011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
100100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
100101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
100110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
100111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
101000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
101001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
101010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
101011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
101100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
101101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
101110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
101111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
110000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
110001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
110010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
110011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
110100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
00
;
6
'b
110101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
110110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
110111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111000
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
01
;
6
'b
111001
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111010
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111011
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111100
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111101
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111110
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
6
'b
111111
:
{
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
}
=
2
'b
10
;
endcase
reg
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
;
always
@
(
CORETSE_AHBlii1I
[
9
:
6
]
)
case
(
{
CORETSE_AHBlii1I
[
9
]
,
CORETSE_AHBlii1I
[
8
]
,
CORETSE_AHBlii1I
[
7
]
,
CORETSE_AHBlii1I
[
6
]
}
)
4
'b
0000
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
01
;
4
'b
0001
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
01
;
4
'b
0010
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
01
;
4
'b
0011
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
10
;
4
'b
0100
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
01
;
4
'b
0101
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
00
;
4
'b
0110
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
00
;
4
'b
0111
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
10
;
4
'b
1000
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
01
;
4
'b
1001
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
00
;
4
'b
1010
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
00
;
4
'b
1011
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
10
;
4
'b
1100
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
01
;
4
'b
1101
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
10
;
4
'b
1110
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
10
;
4
'b
1111
:
{
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
=
2
'b
10
;
endcase
reg
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
;
always
@
(
CORETSE_AHBOloi
or
CORETSE_AHBi0OoI
or
CORETSE_AHBO1OoI
or
CORETSE_AHBI1OoI
or
CORETSE_AHBl1OoI
)
casex
(
{
CORETSE_AHBOloi
,
CORETSE_AHBi0OoI
,
CORETSE_AHBO1OoI
,
CORETSE_AHBI1OoI
,
CORETSE_AHBl1OoI
}
)
5
'b
0_0000
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
00
;
5
'b
1_0000
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
01
;
5
'b
x_1000
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
10
;
5
'b
x_0100
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
00
;
5
'b
x_xx10
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
10
;
5
'b
x_xx01
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
00
;
default
:
{
CORETSE_AHBo1OoI
,
CORETSE_AHBi1OoI
}
=
2
'b
00
;
endcase
assign
CORETSE_AHBO0oi
=
CORETSE_AHBo1OoI
|
CORETSE_AHBi1OoI
;
endmodule
