// REVISION    : $Revision: 1.3 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
petex_top
#
(
parameter
CORETSE_AHBlOI
=
0
)
(
CORETSE_AHBloi0
,
CORETSE_AHBoI
,
CORETSE_AHBOl11
,
CORETSE_AHBOl
,
CORETSE_AHBlO11
,
CORETSE_AHBioO1
,
CORETSE_AHBOiO1
,
CORETSE_AHBIO11
,
CORETSE_AHBIl11
,
CORETSE_AHBll11
,
CORETSE_AHBli01
,
CORETSE_AHBII11
,
CORETSE_AHBol1
)
;
input
CORETSE_AHBloi0
;
input
CORETSE_AHBoI
;
input
[
7
:
0
]
CORETSE_AHBOl11
;
input
CORETSE_AHBOl
;
input
CORETSE_AHBlO11
;
input
[
1
:
0
]
CORETSE_AHBioO1
;
input
[
15
:
0
]
CORETSE_AHBOiO1
;
input
CORETSE_AHBIO11
;
input
CORETSE_AHBIl11
;
input
[
9
:
0
]
CORETSE_AHBll11
;
input
[
2
:
0
]
CORETSE_AHBli01
;
input
CORETSE_AHBII11
;
output
[
9
:
0
]
CORETSE_AHBol1
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBoIlII
;
reg
[
1
:
0
]
CORETSE_AHBiIlII
;
wire
CORETSE_AHBOllII
;
reg
CORETSE_AHBIllII
;
wire
[
7
:
0
]
CORETSE_AHBlllII
;
reg
[
7
:
0
]
CORETSE_AHBollII
;
wire
CORETSE_AHBillII
;
reg
CORETSE_AHBO0lII
;
wire
CORETSE_AHBI0lII
;
reg
CORETSE_AHBl0lII
;
wire
CORETSE_AHBo0lII
;
wire
CORETSE_AHBi0lII
;
wire
CORETSE_AHBO1lII
;
wire
CORETSE_AHBI1lII
;
reg
CORETSE_AHBl1lII
;
wire
CORETSE_AHBo1lII
;
wire
CORETSE_AHBi1lII
;
wire
CORETSE_AHBOolII
;
wire
CORETSE_AHBIolII
;
reg
CORETSE_AHBlolII
;
reg
CORETSE_AHBoolII
;
reg
CORETSE_AHBiolII
;
reg
CORETSE_AHBOilII
;
wire
CORETSE_AHBIilII
;
reg
CORETSE_AHBlilII
;
wire
CORETSE_AHBoilII
;
reg
CORETSE_AHBiilII
;
wire
CORETSE_AHBOO0II
;
reg
CORETSE_AHBIO0II
;
wire
CORETSE_AHBlO0II
;
reg
CORETSE_AHBoO0II
;
wire
CORETSE_AHBiO0II
;
reg
CORETSE_AHBOI0II
;
wire
CORETSE_AHBII0II
;
reg
CORETSE_AHBlI0II
;
wire
CORETSE_AHBoI0II
;
reg
CORETSE_AHBiI0II
;
wire
CORETSE_AHBOl0II
;
wire
CORETSE_AHBIOIOI
;
reg
CORETSE_AHBlOIOI
;
wire
CORETSE_AHBIl0II
;
reg
CORETSE_AHBll0II
;
wire
CORETSE_AHBol0II
;
reg
CORETSE_AHBil0II
;
wire
CORETSE_AHBO00II
;
reg
CORETSE_AHBI00II
;
wire
CORETSE_AHBl00II
;
reg
CORETSE_AHBo00II
;
wire
CORETSE_AHBi00II
;
reg
CORETSE_AHBO10II
;
wire
CORETSE_AHBI10II
;
reg
CORETSE_AHBl10II
;
wire
CORETSE_AHBo10II
;
wire
CORETSE_AHBi10II
;
reg
CORETSE_AHBOo0II
;
wire
CORETSE_AHBIo0II
;
reg
CORETSE_AHBlo0II
;
wire
CORETSE_AHBoo0II
;
reg
CORETSE_AHBio0II
;
wire
[
3
:
0
]
CORETSE_AHBOi0II
;
reg
[
3
:
0
]
CORETSE_AHBIi0II
;
wire
CORETSE_AHBli0II
,
CORETSE_AHBoi0II
;
wire
CORETSE_AHBii0II
;
reg
CORETSE_AHBOO1II
;
wire
[
9
:
0
]
CORETSE_AHBIO1II
;
reg
[
9
:
0
]
CORETSE_AHBlO1II
;
wire
[
7
:
0
]
CORETSE_AHBoO1II
;
reg
[
7
:
0
]
CORETSE_AHBiio
;
wire
[
7
:
0
]
CORETSE_AHBiO1II
;
reg
[
7
:
0
]
CORETSE_AHBOI1II
;
wire
[
9
:
0
]
CORETSE_AHBII1II
;
reg
[
9
:
0
]
CORETSE_AHBlI1II
;
wire
CORETSE_AHBoI1II
;
reg
CORETSE_AHBiI1II
;
wire
[
9
:
0
]
CORETSE_AHBOl1II
;
reg
[
1
:
0
]
CORETSE_AHBIl1II
;
wire
CORETSE_AHBll1II
,
CORETSE_AHBol1II
,
CORETSE_AHBil1II
,
CORETSE_AHBO01II
,
CORETSE_AHBI01II
;
reg
[
15
:
0
]
CORETSE_AHBl01II
;
assign
CORETSE_AHBlllII
=
CORETSE_AHBOl11
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBollII
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
CORETSE_AHBollII
<=
#
CORETSE_AHBIoII
CORETSE_AHBlllII
;
end
assign
CORETSE_AHBillII
=
CORETSE_AHBoI
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBO0lII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO0lII
<=
#
CORETSE_AHBIoII
CORETSE_AHBillII
;
end
assign
CORETSE_AHBI0lII
=
CORETSE_AHBOl
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBl0lII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl0lII
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0lII
;
end
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBoIlII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoIlII
<=
#
CORETSE_AHBIoII
~
CORETSE_AHBoIlII
;
end
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBiIlII
<=
#
CORETSE_AHBIoII
2
'h
3
;
else
CORETSE_AHBiIlII
<=
#
CORETSE_AHBIoII
CORETSE_AHBioO1
;
end
assign
CORETSE_AHBOllII
=
~
CORETSE_AHBIllII
&
(
CORETSE_AHBlOIOI
|
CORETSE_AHBO10II
)
|
CORETSE_AHBIllII
&
~
CORETSE_AHBI00II
&
~
(
~
CORETSE_AHBoIlII
&
CORETSE_AHBil0II
)
&
~
(
~
CORETSE_AHBoIlII
&
CORETSE_AHBlo0II
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBIllII
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBIllII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOllII
;
end
assign
CORETSE_AHBo0lII
=
CORETSE_AHBioO1
==
2
'b
00
;
assign
CORETSE_AHBi0lII
=
CORETSE_AHBioO1
==
2
'b
01
;
assign
CORETSE_AHBO1lII
=
CORETSE_AHBioO1
==
2
'b
10
;
assign
CORETSE_AHBI1lII
=
~
CORETSE_AHBl1lII
&
CORETSE_AHBiIlII
!=
CORETSE_AHBioO1
|
CORETSE_AHBl1lII
&
~
(
(
CORETSE_AHBi1lII
&
~
CORETSE_AHBlolII
)
|
(
CORETSE_AHBOolII
&
~
CORETSE_AHBoolII
)
|
(
CORETSE_AHBIolII
&
~
CORETSE_AHBiolII
)
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBl1lII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1lII
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1lII
;
end
assign
CORETSE_AHBi1lII
=
~
CORETSE_AHBlolII
&
CORETSE_AHBo0lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBlolII
&
~
(
(
~
CORETSE_AHBoolII
&
CORETSE_AHBi0lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
)
|
(
~
CORETSE_AHBiolII
&
CORETSE_AHBO1lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
)
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlolII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlolII
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1lII
;
end
assign
CORETSE_AHBOolII
=
~
CORETSE_AHBoolII
&
CORETSE_AHBi0lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBoolII
&
~
(
(
~
CORETSE_AHBlolII
&
CORETSE_AHBo0lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
)
|
(
~
CORETSE_AHBiolII
&
CORETSE_AHBO1lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
)
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBoolII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoolII
<=
#
CORETSE_AHBIoII
CORETSE_AHBOolII
;
end
assign
CORETSE_AHBIolII
=
~
CORETSE_AHBiolII
&
CORETSE_AHBO1lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBiolII
&
~
(
(
~
CORETSE_AHBlolII
&
CORETSE_AHBo0lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
)
|
(
~
CORETSE_AHBoolII
&
CORETSE_AHBi0lII
&
CORETSE_AHBo1lII
&
CORETSE_AHBl1lII
&
~
CORETSE_AHBoIlII
)
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBiolII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiolII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIolII
;
end
assign
CORETSE_AHBoI1II
=
~
CORETSE_AHBiI1II
&
CORETSE_AHBiolII
&
CORETSE_AHBOolII
|
CORETSE_AHBiI1II
&
~
CORETSE_AHBlilII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBiI1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiI1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI1II
;
end
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBOilII
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBlilII
)
CORETSE_AHBOilII
<=
#
CORETSE_AHBIoII
1
'b
0
;
end
assign
CORETSE_AHBIilII
=
CORETSE_AHBlolII
&
CORETSE_AHBo1lII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBlolII
&
CORETSE_AHBOI0II
|
CORETSE_AHBoolII
&
CORETSE_AHBOilII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBoolII
&
CORETSE_AHBo1lII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBoolII
&
CORETSE_AHBiI0II
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBOilII
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBiI0II
|
CORETSE_AHBiolII
&
CORETSE_AHBI00II
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBiolII
&
CORETSE_AHBo00II
&
~
CORETSE_AHBoIlII
|
CORETSE_AHBiI1II
&
~
CORETSE_AHBoIlII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlilII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlilII
<=
#
CORETSE_AHBIoII
CORETSE_AHBIilII
;
end
assign
CORETSE_AHBoilII
=
CORETSE_AHBlilII
&
~
CORETSE_AHBlI0II
&
CORETSE_AHBlolII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBiilII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiilII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoilII
;
end
assign
CORETSE_AHBOO0II
=
CORETSE_AHBlilII
&
CORETSE_AHBlI0II
&
CORETSE_AHBlolII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBIO0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIO0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBOO0II
;
end
assign
CORETSE_AHBlO0II
=
CORETSE_AHBiilII
|
CORETSE_AHBIO0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBoO0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoO0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBlO0II
;
end
assign
CORETSE_AHBiO0II
=
CORETSE_AHBoO0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBOI0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOI0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO0II
;
end
assign
CORETSE_AHBII0II
=
~
CORETSE_AHBlI0II
&
CORETSE_AHBiilII
|
CORETSE_AHBlI0II
&
~
(
CORETSE_AHBiolII
|
CORETSE_AHBoolII
|
CORETSE_AHBIO0II
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlI0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlI0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBII0II
;
end
assign
CORETSE_AHBoI0II
=
CORETSE_AHBoolII
&
CORETSE_AHBlilII
|
CORETSE_AHBiolII
&
CORETSE_AHBlilII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBiI0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiI0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBoI0II
;
end
assign
CORETSE_AHBOl0II
=
CORETSE_AHBIi0II
==
4
'h
c
&
~
CORETSE_AHBli0II
;
assign
CORETSE_AHBIOIOI
=
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBiI0II
|
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBio0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlOIOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlOIOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOIOI
;
end
assign
CORETSE_AHBIl0II
=
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
CORETSE_AHBlOIOI
|
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
CORETSE_AHBll0II
|
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
CORETSE_AHBl10II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBll0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBll0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl0II
;
end
assign
CORETSE_AHBol0II
=
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBlOIOI
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBll0II
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBl10II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBil0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBil0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0II
;
end
assign
CORETSE_AHBO00II
=
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBil0II
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBlo0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBI00II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI00II
<=
#
CORETSE_AHBIoII
CORETSE_AHBO00II
;
end
assign
CORETSE_AHBl00II
=
CORETSE_AHBiolII
&
CORETSE_AHBI00II
&
~
CORETSE_AHBO0lII
&
CORETSE_AHBoIlII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBo00II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo00II
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00II
;
end
assign
CORETSE_AHBi00II
=
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBiI0II
|
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBio0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBO10II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO10II
<=
#
CORETSE_AHBIoII
CORETSE_AHBi00II
;
end
assign
CORETSE_AHBI10II
=
CORETSE_AHBiolII
&
CORETSE_AHBO10II
|
CORETSE_AHBiolII
&
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBl10II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl10II
<=
#
CORETSE_AHBIoII
CORETSE_AHBI10II
;
end
assign
CORETSE_AHBo10II
=
CORETSE_AHBll0II
&
~
CORETSE_AHBl10II
;
assign
CORETSE_AHBi10II
=
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBlOIOI
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBll0II
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBl10II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBOo0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOo0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBi10II
;
end
assign
CORETSE_AHBIo0II
=
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBOo0II
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
~
CORETSE_AHBl0lII
&
CORETSE_AHBio0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlo0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlo0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo0II
;
end
assign
CORETSE_AHBoo0II
=
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBOo0II
|
CORETSE_AHBiolII
&
~
CORETSE_AHBO0lII
&
CORETSE_AHBl0lII
&
CORETSE_AHBio0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBio0II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBio0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo0II
;
end
assign
CORETSE_AHBiO1II
=
CORETSE_AHBollII
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBOI1II
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
CORETSE_AHBOI1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBiO1II
;
end
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
begin
CORETSE_AHBl01II
<=
#
CORETSE_AHBIoII
16
'h
0
;
end
else
if
(
CORETSE_AHBiilII
)
begin
CORETSE_AHBl01II
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiO1
;
end
else
begin
CORETSE_AHBl01II
<=
#
CORETSE_AHBIoII
CORETSE_AHBl01II
;
end
end
assign
CORETSE_AHBoO1II
=
{
8
{
CORETSE_AHBoO0II
}
}
&
CORETSE_AHBl01II
[
7
:
0
]
|
{
8
{
CORETSE_AHBOI0II
}
}
&
CORETSE_AHBl01II
[
15
:
8
]
|
{
8
{
CORETSE_AHBll0II
}
}
&
CORETSE_AHBOI1II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBiio
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
CORETSE_AHBiio
<=
#
CORETSE_AHBIoII
CORETSE_AHBoO1II
;
end
assign
CORETSE_AHBOi0II
=
{
4
{
CORETSE_AHBiI0II
}
}
&
{
3
'b
000
,
CORETSE_AHBOl0II
}
|
{
4
{
CORETSE_AHBlOIOI
|
CORETSE_AHBO10II
}
}
&
4
'h
8
|
{
4
{
CORETSE_AHBl10II
}
}
&
4
'h
9
|
{
4
{
CORETSE_AHBil0II
|
CORETSE_AHBOo0II
}
}
&
4
'h
a
|
{
4
{
CORETSE_AHBI00II
|
CORETSE_AHBo00II
|
CORETSE_AHBio0II
|
CORETSE_AHBlo0II
}
}
&
4
'h
b
|
{
4
{
CORETSE_AHBlilII
|
CORETSE_AHBOilII
}
}
&
4
'h
c
|
{
4
{
CORETSE_AHBoO0II
|
CORETSE_AHBOI0II
|
CORETSE_AHBo10II
}
}
&
4
'h
d
|
{
4
{
CORETSE_AHBiilII
}
}
&
4
'h
e
|
{
4
{
CORETSE_AHBIO0II
}
}
&
4
'h
f
;
assign
CORETSE_AHBo1lII
=
~
(
CORETSE_AHBlolII
|
CORETSE_AHBoolII
|
CORETSE_AHBiolII
)
|
CORETSE_AHBlolII
&
~
CORETSE_AHBiilII
&
~
CORETSE_AHBIO0II
&
~
CORETSE_AHBoO0II
&
~
CORETSE_AHBOI0II
&
~
CORETSE_AHBlilII
|
CORETSE_AHBlolII
&
CORETSE_AHBOI0II
|
CORETSE_AHBiI0II
|
CORETSE_AHBlOIOI
|
CORETSE_AHBll0II
|
CORETSE_AHBil0II
|
CORETSE_AHBI00II
|
CORETSE_AHBo00II
|
CORETSE_AHBO10II
|
CORETSE_AHBl10II
|
CORETSE_AHBOo0II
|
CORETSE_AHBlo0II
|
CORETSE_AHBio0II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBIi0II
<=
#
CORETSE_AHBIoII
4
'h
c
;
else
CORETSE_AHBIi0II
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi0II
;
end
assign
CORETSE_AHBli0II
=
~
CORETSE_AHBIO11
&
CORETSE_AHBOO1II
;
assign
CORETSE_AHBii0II
=
~
CORETSE_AHBIO11
&
(
CORETSE_AHBOO1II
^
CORETSE_AHBoi0II
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBOO1II
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOO1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBii0II
;
end
t8b10b
CORETSE_AHBo01II
(
.CORETSE_AHBiio
(
CORETSE_AHBiio
)
,
.CORETSE_AHBIi0II
(
CORETSE_AHBIi0II
)
,
.CORETSE_AHBli0II
(
CORETSE_AHBli0II
)
,
.CORETSE_AHBIO1II
(
CORETSE_AHBIO1II
)
,
.CORETSE_AHBoi0II
(
CORETSE_AHBoi0II
)
)
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlO1II
<=
#
CORETSE_AHBIoII
10
'h
0
;
else
CORETSE_AHBlO1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIO1II
;
end
assign
CORETSE_AHBII1II
=
{
10
{
~
CORETSE_AHBlO11
&
~
CORETSE_AHBIl11
}
}
&
CORETSE_AHBlO1II
|
{
10
{
|
CORETSE_AHBli01
&
CORETSE_AHBIl11
}
}
&
CORETSE_AHBOl1II
|
{
10
{
~|
CORETSE_AHBli01
&
CORETSE_AHBIl11
}
}
&
CORETSE_AHBll11
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBlI1II
<=
#
CORETSE_AHBIoII
10
'h
0
;
else
CORETSE_AHBlI1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBII1II
;
end
assign
CORETSE_AHBol1
=
{
10
{
(
CORETSE_AHBlO11
&
~
CORETSE_AHBIl11
)
}
}
&
{
CORETSE_AHBOl
,
CORETSE_AHBoI
,
CORETSE_AHBOl11
[
7
:
0
]
}
|
{
10
{
~
(
CORETSE_AHBlO11
&
~
CORETSE_AHBIl11
)
}
}
&
CORETSE_AHBlI1II
;
always
@
(
posedge
CORETSE_AHBloi0
or
posedge
CORETSE_AHBII11
)
begin
if
(
CORETSE_AHBII11
)
CORETSE_AHBIl1II
<=
#
CORETSE_AHBIoII
2
'h
0
;
else
CORETSE_AHBIl1II
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl1II
+
2
'h
1
;
end
assign
CORETSE_AHBll1II
=
CORETSE_AHBli01
[
2
:
0
]
==
3
'b
001
;
assign
CORETSE_AHBol1II
=
CORETSE_AHBli01
[
2
:
0
]
==
3
'b
010
;
assign
CORETSE_AHBil1II
=
CORETSE_AHBli01
[
2
:
0
]
==
3
'b
011
;
assign
CORETSE_AHBO01II
=
CORETSE_AHBli01
[
2
:
0
]
==
3
'b
100
;
assign
CORETSE_AHBI01II
=
CORETSE_AHBli01
[
2
:
0
]
==
3
'b
101
;
assign
CORETSE_AHBOl1II
=
{
10
{
(
CORETSE_AHBll1II
)
}
}
&
10
'h
255
|
{
10
{
(
CORETSE_AHBol1II
&
~
CORETSE_AHBIl1II
[
0
]
)
}
}
&
10
'h
17c
|
{
10
{
(
CORETSE_AHBol1II
&
CORETSE_AHBIl1II
[
0
]
)
}
}
&
10
'h
283
|
{
10
{
(
CORETSE_AHBil1II
)
}
}
&
10
'h
3e0
|
{
10
{
(
CORETSE_AHBO01II
&
CORETSE_AHBIl1II
==
2
'h
0
)
}
}
&
10
'h
17c
|
{
10
{
(
CORETSE_AHBO01II
&
CORETSE_AHBIl1II
==
2
'h
1
)
}
}
&
10
'h
0c9
|
{
10
{
(
CORETSE_AHBO01II
&
CORETSE_AHBIl1II
==
2
'h
2
)
}
}
&
10
'h
0e5
|
{
10
{
(
CORETSE_AHBO01II
&
CORETSE_AHBIl1II
==
2
'h
3
)
}
}
&
10
'h
2a3
|
{
10
{
(
CORETSE_AHBI01II
)
}
}
&
10
'h
07c
;
endmodule
