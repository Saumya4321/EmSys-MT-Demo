// REVISION    : $Revision: 1.4 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_core
#
(
parameter
CORETSE_AHBlOI
=
1
'b
0
,
parameter
MDIO_PHYID
=
18
)
(
CORETSE_AHBIi0
,
CORETSE_AHBli0
,
CORETSE_AHBoi0
,
CORETSE_AHBii0
,
CORETSE_AHBlO1
,
CORETSE_AHBiO1
,
CORETSE_AHBII
,
CORETSE_AHBoI
,
CORETSE_AHBOl
,
CORETSE_AHBo11
,
CORETSE_AHBi01
,
CORETSE_AHBO11
,
CORETSE_AHBI11
,
CORETSE_AHBl11
,
CORETSE_AHBll1
,
CORETSE_AHBil1
,
CORETSE_AHBl01
,
CORETSE_AHBOI1
,
CORETSE_AHBII1
,
CORETSE_AHBOO1
,
CORETSE_AHBIO1
,
CORETSE_AHBlI1
,
CORETSE_AHBoI1
,
CORETSE_AHBiI1
,
CORETSE_AHBOl1
,
CORETSE_AHBol1
,
CORETSE_AHBIl1
,
CORETSE_AHBlI
,
CORETSE_AHBiI
,
CORETSE_AHBIl
,
CORETSE_AHBO01
,
CORETSE_AHBol
,
CORETSE_AHBo01
,
CORETSE_AHBI01
,
CORETSE_AHBoO1
,
CORETSE_AHBi11
,
CORETSE_AHBOo1
)
;
input
CORETSE_AHBIi0
;
input
CORETSE_AHBli0
;
input
CORETSE_AHBoi0
;
input
CORETSE_AHBii0
;
input
CORETSE_AHBlO1
;
input
CORETSE_AHBiO1
;
input
[
7
:
0
]
CORETSE_AHBII
;
input
CORETSE_AHBoI
;
input
CORETSE_AHBOl
;
input
[
1
:
0
]
CORETSE_AHBo11
;
input
CORETSE_AHBi01
;
input
CORETSE_AHBO11
;
input
CORETSE_AHBI11
;
input
CORETSE_AHBl11
;
input
CORETSE_AHBll1
;
input
[
9
:
0
]
CORETSE_AHBil1
;
input
CORETSE_AHBOI1
;
input
CORETSE_AHBII1
;
input
CORETSE_AHBOO1
;
input
CORETSE_AHBIO1
;
input
CORETSE_AHBl01
;
output
CORETSE_AHBlI1
;
output
CORETSE_AHBoI1
;
output
CORETSE_AHBiI1
;
output
CORETSE_AHBOl1
;
output
[
9
:
0
]
CORETSE_AHBol1
;
output
CORETSE_AHBIl1
;
output
[
7
:
0
]
CORETSE_AHBlI
;
output
CORETSE_AHBiI
;
output
CORETSE_AHBIl
;
output
CORETSE_AHBO01
;
output
CORETSE_AHBol
;
output
CORETSE_AHBo01
;
output
CORETSE_AHBI01
;
output
CORETSE_AHBoO1
;
output
reg
[
9
:
0
]
CORETSE_AHBi11
;
output
CORETSE_AHBOo1
;
wire
[
7
:
0
]
CORETSE_AHBloo0
;
wire
CORETSE_AHBooo0
;
wire
CORETSE_AHBioo0
;
wire
[
7
:
0
]
CORETSE_AHBI0i0
;
wire
CORETSE_AHBo110
;
wire
CORETSE_AHBl0i0
;
wire
[
15
:
0
]
CORETSE_AHBO110
;
wire
[
1
:
0
]
CORETSE_AHBI110
;
wire
[
1
:
0
]
CORETSE_AHBl110
;
wire
[
7
:
0
]
CORETSE_AHBOo10
;
wire
CORETSE_AHBIo10
;
wire
CORETSE_AHBlo10
;
wire
[
2
:
0
]
CORETSE_AHBIoo0
;
wire
[
3
:
0
]
CORETSE_AHBi110
;
wire
[
2
:
0
]
CORETSE_AHBIio0
;
wire
[
3
:
0
]
CORETSE_AHBio10
;
wire
CORETSE_AHBOio0
;
wire
CORETSE_AHBoo10
;
wire
CORETSE_AHBi010
;
wire
CORETSE_AHBoO10
;
wire
CORETSE_AHBiO10
;
wire
CORETSE_AHBOI10
;
wire
[
8
:
0
]
CORETSE_AHBI1i0
;
wire
CORETSE_AHBl1i0
;
always
@
(
posedge
CORETSE_AHBli0
or
posedge
CORETSE_AHBIi0
)
begin
if
(
CORETSE_AHBIi0
==
1
'b
1
)
CORETSE_AHBi11
<=
10
'h
0
;
else
CORETSE_AHBi11
<=
{
CORETSE_AHBl1i0
,
CORETSE_AHBI1i0
[
8
:
0
]
}
;
end
msgmii_clkrst
CORETSE_AHBo1i0
(
.CORETSE_AHBIi0
(
CORETSE_AHBIi0
)
,
.CORETSE_AHBll1
(
CORETSE_AHBll1
)
,
.CORETSE_AHBli0
(
CORETSE_AHBli0
)
,
.CORETSE_AHBoi0
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBii0
(
CORETSE_AHBii0
)
,
.CORETSE_AHBlO1
(
CORETSE_AHBlO1
)
,
.CORETSE_AHBiO1
(
CORETSE_AHBiO1
)
,
.CORETSE_AHBoO10
(
CORETSE_AHBoO10
)
,
.CORETSE_AHBiO10
(
CORETSE_AHBiO10
)
,
.CORETSE_AHBOI10
(
CORETSE_AHBOI10
)
,
.CORETSE_AHBlI1
(
CORETSE_AHBlI1
)
,
.CORETSE_AHBoI1
(
CORETSE_AHBoI1
)
,
.CORETSE_AHBoO1
(
CORETSE_AHBoO1
)
)
;
msgmii_cnvtxi
CORETSE_AHBi1i0
(
.CORETSE_AHBiO10
(
CORETSE_AHBiO10
)
,
.CORETSE_AHBoi0
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBo11
(
CORETSE_AHBo11
)
,
.CORETSE_AHBII
(
CORETSE_AHBII
)
,
.CORETSE_AHBoI
(
CORETSE_AHBoI
)
,
.CORETSE_AHBOl
(
CORETSE_AHBOl
)
,
.CORETSE_AHBIoo0
(
CORETSE_AHBIoo0
)
,
.CORETSE_AHBloo0
(
CORETSE_AHBloo0
)
,
.CORETSE_AHBooo0
(
CORETSE_AHBooo0
)
,
.CORETSE_AHBioo0
(
CORETSE_AHBioo0
)
,
.CORETSE_AHBOio0
(
CORETSE_AHBOio0
)
,
.CORETSE_AHBIio0
(
CORETSE_AHBIio0
)
)
;
msgmii_cnvtxo
CORETSE_AHBOoi0
(
.CORETSE_AHBoO10
(
CORETSE_AHBoO10
)
,
.CORETSE_AHBli0
(
CORETSE_AHBli0
)
,
.CORETSE_AHBo11
(
CORETSE_AHBo11
)
,
.CORETSE_AHBloo0
(
CORETSE_AHBloo0
)
,
.CORETSE_AHBooo0
(
CORETSE_AHBooo0
)
,
.CORETSE_AHBioo0
(
CORETSE_AHBioo0
)
,
.CORETSE_AHBOio0
(
CORETSE_AHBOio0
)
,
.CORETSE_AHBIio0
(
CORETSE_AHBIio0
)
,
.CORETSE_AHBIoo0
(
CORETSE_AHBIoo0
)
,
.CORETSE_AHBI0i0
(
CORETSE_AHBI0i0
)
,
.CORETSE_AHBo110
(
CORETSE_AHBo110
)
,
.CORETSE_AHBl0i0
(
CORETSE_AHBl0i0
)
,
.CORETSE_AHBIl1
(
CORETSE_AHBIl1
)
)
;
msgmii_tbi
#
(
.CORETSE_AHBlOI
(
CORETSE_AHBlOI
)
)
CORETSE_AHBIoi0
(
.CORETSE_AHBloi0
(
CORETSE_AHBli0
)
,
.CORETSE_AHBII
(
CORETSE_AHBI0i0
)
,
.CORETSE_AHBoI
(
CORETSE_AHBo110
)
,
.CORETSE_AHBOl
(
CORETSE_AHBl0i0
)
,
.CORETSE_AHBII1
(
CORETSE_AHBII1
)
,
.CORETSE_AHBOI1
(
CORETSE_AHBOI1
)
,
.CORETSE_AHBIO1
(
CORETSE_AHBIO1
)
,
.CORETSE_AHBOO1
(
CORETSE_AHBOO1
)
,
.CORETSE_AHBil1
(
CORETSE_AHBil1
)
,
.CORETSE_AHBl01
(
CORETSE_AHBl01
)
,
.CORETSE_AHBi01
(
CORETSE_AHBi01
)
,
.CORETSE_AHBO11
(
CORETSE_AHBO11
)
,
.CORETSE_AHBI11
(
CORETSE_AHBI11
)
,
.CORETSE_AHBl11
(
CORETSE_AHBl11
)
,
.CORETSE_AHBooi0
(
MDIO_PHYID
[
4
:
0
]
)
,
.CORETSE_AHBioi0
(
CORETSE_AHBIi0
)
,
.CORETSE_AHBll1
(
CORETSE_AHBll1
)
,
.CORETSE_AHBol1
(
CORETSE_AHBol1
)
,
.CORETSE_AHBOl1
(
CORETSE_AHBOl1
)
,
.CORETSE_AHBiI1
(
CORETSE_AHBiI1
)
,
.CORETSE_AHBi010
(
CORETSE_AHBi010
)
,
.CORETSE_AHBOii0
(
CORETSE_AHBO110
)
,
.CORETSE_AHBIii0
(
CORETSE_AHBI110
)
,
.CORETSE_AHBlii0
(
CORETSE_AHBl110
)
,
.CORETSE_AHBo01
(
CORETSE_AHBo01
)
,
.CORETSE_AHBoii0
(
)
,
.CORETSE_AHBiii0
(
CORETSE_AHBI01
)
,
.CORETSE_AHBOOO1
(
)
,
.CORETSE_AHBIOO1
(
CORETSE_AHBOo1
)
,
.CORETSE_AHBl1i0
(
CORETSE_AHBl1i0
)
,
.CORETSE_AHBI1i0
(
CORETSE_AHBI1i0
)
)
;
msgmii_cnvrxi
CORETSE_AHBlOO1
(
.CORETSE_AHBi010
(
CORETSE_AHBi010
)
,
.CORETSE_AHBOO1
(
CORETSE_AHBOO1
)
,
.CORETSE_AHBo11
(
CORETSE_AHBo11
)
,
.CORETSE_AHBO110
(
CORETSE_AHBO110
)
,
.CORETSE_AHBI110
(
CORETSE_AHBI110
)
,
.CORETSE_AHBl110
(
CORETSE_AHBl110
)
,
.CORETSE_AHBo110
(
CORETSE_AHBo110
)
,
.CORETSE_AHBi110
(
CORETSE_AHBi110
)
,
.CORETSE_AHBOo10
(
CORETSE_AHBOo10
)
,
.CORETSE_AHBIo10
(
CORETSE_AHBIo10
)
,
.CORETSE_AHBlo10
(
CORETSE_AHBlo10
)
,
.CORETSE_AHBO01
(
CORETSE_AHBO01
)
,
.CORETSE_AHBol
(
CORETSE_AHBol
)
,
.CORETSE_AHBoo10
(
CORETSE_AHBoo10
)
,
.CORETSE_AHBio10
(
CORETSE_AHBio10
)
)
;
msgmii_cnvrxo
CORETSE_AHBoOO1
(
.CORETSE_AHBOI10
(
CORETSE_AHBOI10
)
,
.CORETSE_AHBii0
(
CORETSE_AHBii0
)
,
.CORETSE_AHBo11
(
CORETSE_AHBo11
)
,
.CORETSE_AHBOo10
(
CORETSE_AHBOo10
)
,
.CORETSE_AHBIo10
(
CORETSE_AHBIo10
)
,
.CORETSE_AHBlo10
(
CORETSE_AHBlo10
)
,
.CORETSE_AHBoo10
(
CORETSE_AHBoo10
)
,
.CORETSE_AHBio10
(
CORETSE_AHBio10
)
,
.CORETSE_AHBlI
(
CORETSE_AHBlI
)
,
.CORETSE_AHBiI
(
CORETSE_AHBiI
)
,
.CORETSE_AHBIl
(
CORETSE_AHBIl
)
,
.CORETSE_AHBi110
(
CORETSE_AHBi110
)
)
;
endmodule
