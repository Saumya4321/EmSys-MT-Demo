// REVISION    : $Revision: 1.7 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
permc_top
(
CORETSE_AHBo111
,
CORETSE_AHBi1Oo
,
CORETSE_AHBI1Io
,
CORETSE_AHBl1Io
,
CORETSE_AHBo1Io
,
CORETSE_AHBi1Io
,
CORETSE_AHBOoIo
,
CORETSE_AHBIoIo
,
CORETSE_AHBoo01
,
CORETSE_AHBOli1
,
CORETSE_AHBiIi1
,
CORETSE_AHBll00
,
CORETSE_AHBIli1
,
CORETSE_AHBi0Oo
,
CORETSE_AHBO0Io
,
CORETSE_AHBOiIo
,
CORETSE_AHBo0o
,
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
,
CORETSE_AHBo1o
,
CORETSE_AHBl1o
,
CORETSE_AHBIiIo
,
CORETSE_AHBliIo
,
CORETSE_AHBoiIo
,
CORETSE_AHBIl00
)
;
input
CORETSE_AHBo111
,
CORETSE_AHBi1Oo
;
input
[
7
:
0
]
CORETSE_AHBI1Io
;
input
CORETSE_AHBl1Io
,
CORETSE_AHBo1Io
,
CORETSE_AHBi1Io
;
input
CORETSE_AHBOoIo
;
input
[
32
:
0
]
CORETSE_AHBIoIo
;
input
[
1
:
0
]
CORETSE_AHBoo01
;
input
CORETSE_AHBiIi1
;
input
[
47
:
0
]
CORETSE_AHBll00
;
input
CORETSE_AHBIli1
;
input
CORETSE_AHBi0Oo
;
input
CORETSE_AHBO0Io
;
input
CORETSE_AHBOli1
;
output
[
7
:
0
]
CORETSE_AHBo0o
;
output
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
;
output
CORETSE_AHBo1o
;
output
[
32
:
0
]
CORETSE_AHBl1o
;
output
CORETSE_AHBOiIo
;
output
CORETSE_AHBIiIo
,
CORETSE_AHBliIo
,
CORETSE_AHBoiIo
,
CORETSE_AHBIl00
;
reg
[
7
:
0
]
CORETSE_AHBo0o
;
reg
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
;
reg
CORETSE_AHBo1o
;
reg
[
32
:
0
]
CORETSE_AHBl1o
;
reg
CORETSE_AHBOiIo
;
reg
CORETSE_AHBIiIo
,
CORETSE_AHBliIo
,
CORETSE_AHBoiIo
,
CORETSE_AHBIl00
;
parameter
CORETSE_AHBIoII
=
1
;
wire
[
4
:
0
]
CORETSE_AHBOooOI
;
wire
CORETSE_AHBIooOI
,
CORETSE_AHBlooOI
;
wire
[
4
:
0
]
CORETSE_AHBoooOI
;
reg
[
4
:
0
]
CORETSE_AHBiooOI
;
wire
CORETSE_AHBOioOI
,
CORETSE_AHBIioOI
,
CORETSE_AHBlioOI
,
CORETSE_AHBoioOI
;
wire
CORETSE_AHBiioOI
,
CORETSE_AHBOOiOI
,
CORETSE_AHBIOiOI
;
wire
CORETSE_AHBlOiOI
,
CORETSE_AHBoOiOI
,
CORETSE_AHBiOiOI
,
CORETSE_AHBOIiOI
;
wire
CORETSE_AHBIIiOI
,
CORETSE_AHBlIiOI
;
wire
CORETSE_AHBoIiOI
,
CORETSE_AHBiIiOI
,
CORETSE_AHBOliOI
,
CORETSE_AHBIliOI
;
wire
CORETSE_AHBlliOI
,
CORETSE_AHBoliOI
;
wire
CORETSE_AHBiliOI
,
CORETSE_AHBO0iOI
,
CORETSE_AHBI0iOI
,
CORETSE_AHBl0iOI
;
wire
CORETSE_AHBo0iOI
,
CORETSE_AHBi0iOI
;
wire
CORETSE_AHBO1iOI
,
CORETSE_AHBI1iOI
;
wire
CORETSE_AHBIo1OI
;
reg
CORETSE_AHBOl00
;
wire
CORETSE_AHBl1iOI
;
wire
CORETSE_AHBo1iOI
;
reg
CORETSE_AHBi1iOI
;
wire
[
15
:
0
]
CORETSE_AHBOoiOI
;
reg
[
15
:
0
]
CORETSE_AHBIoiOI
;
wire
CORETSE_AHBloiOI
;
wire
[
15
:
0
]
CORETSE_AHBooiOI
;
reg
[
15
:
0
]
CORETSE_AHBioiOI
;
wire
CORETSE_AHBOiiOI
;
reg
CORETSE_AHBIiiOI
;
wire
CORETSE_AHBliiOI
,
CORETSE_AHBoiiOI
;
reg
CORETSE_AHBiiiOI
,
CORETSE_AHBOOOII
;
wire
[
15
:
0
]
CORETSE_AHBIOOII
;
reg
[
15
:
0
]
CORETSE_AHBlOOII
;
wire
CORETSE_AHBoOOII
,
CORETSE_AHBiOOII
;
wire
[
6
:
0
]
CORETSE_AHBOIOII
;
reg
[
6
:
0
]
CORETSE_AHBIIOII
;
wire
CORETSE_AHBlIOII
;
reg
CORETSE_AHBoIOII
;
wire
CORETSE_AHBiIOII
,
CORETSE_AHBOlOII
,
CORETSE_AHBIlOII
;
reg
CORETSE_AHBllOII
;
reg
CORETSE_AHBolOII
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
begin
CORETSE_AHBllOII
<=
#
CORETSE_AHBIoII
1
'h
0
;
CORETSE_AHBolOII
<=
#
CORETSE_AHBIoII
1
'h
0
;
end
else
begin
CORETSE_AHBllOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0Io
;
CORETSE_AHBolOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBllOII
;
end
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBo0o
[
7
:
0
]
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBo0o
[
7
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1Io
[
7
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBi0o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBi0o
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1Io
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBO1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBO1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1Io
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBI1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBI1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1Io
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBo1o
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBo1o
<=
#
CORETSE_AHBIoII
CORETSE_AHBOoIo
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBl1o
[
32
:
0
]
<=
#
CORETSE_AHBIoII
33
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBl1o
[
32
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoIo
[
32
:
0
]
;
end
assign
CORETSE_AHBOooOI
[
4
:
0
]
=
5
'b
0_0000
;
assign
CORETSE_AHBIooOI
=
CORETSE_AHBOoIo
;
assign
CORETSE_AHBlooOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
!=
5
'b
1_0010
;
assign
CORETSE_AHBoooOI
[
4
:
0
]
=
{
5
{
CORETSE_AHBIooOI
}
}
&
CORETSE_AHBOooOI
[
4
:
0
]
|
{
5
{
~
CORETSE_AHBIooOI
&
CORETSE_AHBlooOI
}
}
&
CORETSE_AHBiooOI
[
4
:
0
]
+
1
'b
1
|
{
5
{
~
CORETSE_AHBIooOI
&
~
CORETSE_AHBlooOI
}
}
&
CORETSE_AHBiooOI
[
4
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBiooOI
[
4
:
0
]
<=
#
CORETSE_AHBIoII
5
'b
0_0000
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiooOI
[
4
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBoooOI
[
4
:
0
]
;
end
assign
CORETSE_AHBOioOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_0000
;
assign
CORETSE_AHBIioOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_0001
;
assign
CORETSE_AHBlioOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_0010
;
assign
CORETSE_AHBoioOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_0011
;
assign
CORETSE_AHBiioOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_0100
;
assign
CORETSE_AHBOOiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_0101
;
assign
CORETSE_AHBIOiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
>
5
'b
0_0101
;
assign
CORETSE_AHBlOiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_1100
;
assign
CORETSE_AHBoOiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_1101
;
assign
CORETSE_AHBiOiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_1110
;
assign
CORETSE_AHBOIiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
0_1111
;
assign
CORETSE_AHBIIiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
1_0000
;
assign
CORETSE_AHBlIiOI
=
CORETSE_AHBl1Io
&
CORETSE_AHBiooOI
[
4
:
0
]
==
5
'b
1_0001
;
assign
CORETSE_AHBoIiOI
=
CORETSE_AHBOioOI
&
(
8
'h
01
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBiIiOI
=
CORETSE_AHBIioOI
&
(
8
'h
80
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBOliOI
=
CORETSE_AHBlioOI
&
(
8
'h
c2
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBIliOI
=
CORETSE_AHBoioOI
&
(
8
'h
00
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBlliOI
=
CORETSE_AHBiioOI
&
(
8
'h
00
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBoliOI
=
CORETSE_AHBOOiOI
&
(
8
'h
01
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBiliOI
=
CORETSE_AHBOioOI
&
(
CORETSE_AHBll00
[
47
:
40
]
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBO0iOI
=
CORETSE_AHBIioOI
&
(
CORETSE_AHBll00
[
39
:
32
]
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBI0iOI
=
CORETSE_AHBlioOI
&
(
CORETSE_AHBll00
[
31
:
24
]
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBl0iOI
=
CORETSE_AHBoioOI
&
(
CORETSE_AHBll00
[
23
:
16
]
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBo0iOI
=
CORETSE_AHBiioOI
&
(
CORETSE_AHBll00
[
15
:
8
]
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBi0iOI
=
CORETSE_AHBOOiOI
&
(
CORETSE_AHBll00
[
7
:
0
]
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBO1iOI
=
CORETSE_AHBlOiOI
&
(
8
'h
88
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBI1iOI
=
CORETSE_AHBoOiOI
&
(
8
'h
08
==
CORETSE_AHBI1Io
[
7
:
0
]
)
;
assign
CORETSE_AHBIo1OI
=
~
CORETSE_AHBOl00
&
CORETSE_AHBOioOI
&
CORETSE_AHBoIiOI
|
CORETSE_AHBOl00
&
CORETSE_AHBOioOI
&
CORETSE_AHBoIiOI
|
CORETSE_AHBOl00
&
CORETSE_AHBIioOI
&
CORETSE_AHBiIiOI
|
CORETSE_AHBOl00
&
CORETSE_AHBlioOI
&
CORETSE_AHBOliOI
|
CORETSE_AHBOl00
&
CORETSE_AHBoioOI
&
CORETSE_AHBIliOI
|
CORETSE_AHBOl00
&
CORETSE_AHBiioOI
&
CORETSE_AHBlliOI
|
CORETSE_AHBOl00
&
CORETSE_AHBOOiOI
&
CORETSE_AHBoliOI
|
CORETSE_AHBOl00
&
(
CORETSE_AHBIOiOI
|
~
CORETSE_AHBl1Io
)
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBOl00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOl00
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo1OI
;
end
assign
CORETSE_AHBl1iOI
=
~
CORETSE_AHBIl00
&
CORETSE_AHBOioOI
&
CORETSE_AHBiliOI
|
CORETSE_AHBIl00
&
CORETSE_AHBIioOI
&
CORETSE_AHBO0iOI
|
CORETSE_AHBIl00
&
CORETSE_AHBlioOI
&
CORETSE_AHBI0iOI
|
CORETSE_AHBIl00
&
CORETSE_AHBoioOI
&
CORETSE_AHBl0iOI
|
CORETSE_AHBIl00
&
CORETSE_AHBiioOI
&
CORETSE_AHBo0iOI
|
CORETSE_AHBIl00
&
CORETSE_AHBOOiOI
&
CORETSE_AHBi0iOI
|
CORETSE_AHBIl00
&
CORETSE_AHBIOiOI
|
CORETSE_AHBIl00
&
~
CORETSE_AHBl1Io
&
~
CORETSE_AHBo1o
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBIl00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIl00
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1iOI
;
end
assign
CORETSE_AHBo1iOI
=
~
CORETSE_AHBi1iOI
&
CORETSE_AHBlOiOI
&
CORETSE_AHBO1iOI
|
CORETSE_AHBi1iOI
&
CORETSE_AHBoOiOI
&
CORETSE_AHBI1iOI
|
CORETSE_AHBi1iOI
&
~
(
CORETSE_AHBlOiOI
&
~
CORETSE_AHBO1iOI
|
CORETSE_AHBoOiOI
&
~
CORETSE_AHBI1iOI
)
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBi1iOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBi1iOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1iOI
;
end
assign
CORETSE_AHBOoiOI
[
15
:
0
]
=
{
16
{
CORETSE_AHBiOiOI
}
}
&
{
CORETSE_AHBI1Io
[
7
:
0
]
,
CORETSE_AHBIoiOI
[
7
:
0
]
}
|
{
16
{
CORETSE_AHBOIiOI
}
}
&
{
CORETSE_AHBIoiOI
[
15
:
8
]
,
CORETSE_AHBI1Io
[
7
:
0
]
}
|
{
16
{
~
CORETSE_AHBiOiOI
&
~
CORETSE_AHBOIiOI
}
}
&
{
CORETSE_AHBIoiOI
[
15
:
8
]
,
CORETSE_AHBIoiOI
[
7
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBIoiOI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIoiOI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOoiOI
[
15
:
0
]
;
end
assign
CORETSE_AHBloiOI
=
CORETSE_AHBIoiOI
[
15
:
0
]
==
16
'h
0001
;
assign
CORETSE_AHBooiOI
[
15
:
0
]
=
{
16
{
CORETSE_AHBIIiOI
}
}
&
{
CORETSE_AHBI1Io
[
7
:
0
]
,
CORETSE_AHBioiOI
[
7
:
0
]
}
|
{
16
{
CORETSE_AHBlIiOI
}
}
&
{
CORETSE_AHBioiOI
[
15
:
8
]
,
CORETSE_AHBI1Io
[
7
:
0
]
}
|
{
16
{
~
CORETSE_AHBIIiOI
&
~
CORETSE_AHBlIiOI
}
}
&
{
CORETSE_AHBioiOI
[
15
:
8
]
,
CORETSE_AHBioiOI
[
7
:
0
]
}
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBioiOI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBioiOI
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBooiOI
[
15
:
0
]
;
end
assign
CORETSE_AHBOiiOI
=
(
CORETSE_AHBOl00
|
CORETSE_AHBIl00
)
&
CORETSE_AHBi1iOI
&
CORETSE_AHBloiOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBIiiOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIiiOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiiOI
;
end
assign
CORETSE_AHBliiOI
=
CORETSE_AHBIiiOI
&
CORETSE_AHBOoIo
&
CORETSE_AHBIoIo
[
23
]
&
CORETSE_AHBIoIo
[
15
:
0
]
>=
16
'h
0040
&
CORETSE_AHBIoIo
[
15
:
0
]
<=
16
'h
5dc
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBiiiOI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBiiiOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBliiOI
;
end
assign
CORETSE_AHBoiiOI
=
CORETSE_AHBlIOII
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBOOOII
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOOOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiiOI
;
end
assign
CORETSE_AHBIOOII
[
15
:
0
]
=
{
16
{
CORETSE_AHBiiiOI
}
}
&
CORETSE_AHBioiOI
[
15
:
0
]
|
{
16
{
~
CORETSE_AHBiiiOI
&
CORETSE_AHBOOOII
&
|
CORETSE_AHBlOOII
}
}
&
CORETSE_AHBlOOII
[
15
:
0
]
-
1
'b
1
|
{
16
{
~
CORETSE_AHBiiiOI
&
~
CORETSE_AHBOOOII
}
}
&
CORETSE_AHBlOOII
[
15
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBlOOII
[
15
:
0
]
<=
#
CORETSE_AHBIoII
16
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBlOOII
[
15
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOOII
[
15
:
0
]
;
end
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBOiIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBOiIo
<=
#
CORETSE_AHBIoII
|
CORETSE_AHBlOOII
[
15
:
0
]
&
CORETSE_AHBiIi1
|
CORETSE_AHBOli1
;
end
assign
CORETSE_AHBoOOII
=
CORETSE_AHBiiiOI
|
CORETSE_AHBoIOII
;
assign
CORETSE_AHBiOOII
=
|
CORETSE_AHBlOOII
[
15
:
0
]
;
assign
CORETSE_AHBOIOII
[
6
:
0
]
=
{
7
{
~
CORETSE_AHBoOOII
&
CORETSE_AHBiOOII
&
CORETSE_AHBolOII
}
}
&
CORETSE_AHBIIOII
[
6
:
0
]
+
1
'b
1
|
{
7
{
~
CORETSE_AHBoOOII
&
CORETSE_AHBiOOII
&
~
CORETSE_AHBolOII
}
}
&
CORETSE_AHBIIOII
[
6
:
0
]
|
{
7
{
~
CORETSE_AHBoOOII
&
~
CORETSE_AHBiOOII
}
}
&
CORETSE_AHBIIOII
[
6
:
0
]
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBIIOII
[
6
:
0
]
<=
#
CORETSE_AHBIoII
7
'h
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIIOII
[
6
:
0
]
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIOII
[
6
:
0
]
;
end
assign
CORETSE_AHBlIOII
=
~
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBIIOII
[
6
:
0
]
==
7
'h
7e
&
CORETSE_AHBiOOII
&
CORETSE_AHBolOII
|
CORETSE_AHBoo01
[
1
]
&
CORETSE_AHBIIOII
[
6
:
0
]
==
7
'h
3e
&
CORETSE_AHBiOOII
&
CORETSE_AHBolOII
|
CORETSE_AHBIli1
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBoIOII
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoIOII
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIOII
;
end
assign
CORETSE_AHBiIOII
=
CORETSE_AHBi1iOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBIiIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBIiIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIOII
;
end
assign
CORETSE_AHBOlOII
=
(
CORETSE_AHBOl00
|
CORETSE_AHBIl00
)
&
CORETSE_AHBi1iOI
&
CORETSE_AHBloiOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBliIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBliIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOlOII
;
end
assign
CORETSE_AHBIlOII
=
CORETSE_AHBi1iOI
&
~
CORETSE_AHBloiOI
;
always
@
(
posedge
CORETSE_AHBo111
or
posedge
CORETSE_AHBi0Oo
)
begin
if
(
CORETSE_AHBi0Oo
)
CORETSE_AHBoiIo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBi1Oo
)
CORETSE_AHBoiIo
<=
#
CORETSE_AHBIoII
CORETSE_AHBIlOII
;
end
endmodule
