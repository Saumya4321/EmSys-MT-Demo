// REVISION    : $Revision: 1.8 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
amcxtfif_sys
#
(
parameter
TABITS
=
12
,
parameter
CORETSE_AHBIo1
=
32
,
parameter
CORETSE_AHBlo1
=
$clog2
(
CORETSE_AHBIo1
/
8
)
,
parameter
CORETSE_AHBoOI
=
0
)
(
CORETSE_AHBoi0
,
CORETSE_AHBllo
,
CORETSE_AHBO0II
,
CORETSE_AHBOOII
,
CORETSE_AHBili
,
CORETSE_AHBolo
,
CORETSE_AHBilo
,
CORETSE_AHBO0o
,
CORETSE_AHBI0o
,
CORETSE_AHBOoi
,
CORETSE_AHBIoi
,
CORETSE_AHBloi
,
CORETSE_AHBlIII
,
CORETSE_AHBoIII
,
CORETSE_AHBiOOI
,
CORETSE_AHBoli
,
CORETSE_AHBiio
,
CORETSE_AHBOOi
,
CORETSE_AHBIOi
,
CORETSE_AHBlOi
,
CORETSE_AHBoOi
,
CORETSE_AHBiOi
,
CORETSE_AHBOIi
,
CORETSE_AHBIIi
,
CORETSE_AHBl1i
,
CORETSE_AHBo1i
,
CORETSE_AHBi1i
,
CORETSE_AHBIlOI
,
CORETSE_AHBllOI
)
;
input
CORETSE_AHBoi0
;
input
CORETSE_AHBllo
;
input
CORETSE_AHBO0II
;
input
CORETSE_AHBOOII
;
input
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBili
;
input
CORETSE_AHBolo
;
input
CORETSE_AHBilo
;
input
CORETSE_AHBO0o
;
input
CORETSE_AHBI0o
;
input
[
TABITS
:
0
]
CORETSE_AHBOoi
;
input
CORETSE_AHBIoi
;
input
CORETSE_AHBloi
;
input
[
TABITS
+
1
:
0
]
CORETSE_AHBlIII
;
input
CORETSE_AHBoIII
;
output
CORETSE_AHBiOOI
;
output
[
(
TABITS
-
1
)
:
0
]
CORETSE_AHBoli
;
output
[
7
:
0
]
CORETSE_AHBiio
;
output
CORETSE_AHBOOi
;
output
CORETSE_AHBIOi
;
output
CORETSE_AHBlOi
;
output
CORETSE_AHBoOi
;
output
CORETSE_AHBiOi
;
output
CORETSE_AHBOIi
;
output
CORETSE_AHBIIi
;
output
CORETSE_AHBl1i
;
output
[
TABITS
:
0
]
CORETSE_AHBo1i
;
output
CORETSE_AHBi1i
;
output
CORETSE_AHBIlOI
;
output
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBllOI
;
parameter
CORETSE_AHBol0I
=
{
(
TABITS
+
1
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBiOiI
=
{
(
TABITS
+
(
CORETSE_AHBlo1
+
1
)
)
{
1
'b
0
}
}
;
parameter
CORETSE_AHBIoII
=
1
;
reg
[
5
:
0
]
CORETSE_AHBOIiI
;
reg
CORETSE_AHBIIiI
;
wire
CORETSE_AHBlIiI
;
reg
CORETSE_AHBoIiI
;
reg
CORETSE_AHBiIiI
;
reg
CORETSE_AHBOliI
;
reg
[
TABITS
:
0
]
CORETSE_AHBIliI
;
wire
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBl00I
;
wire
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBlliI
;
wire
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBoliI
;
wire
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBo00I
;
reg
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBiliI
;
reg
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBO0iI
;
reg
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBI0iI
;
reg
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBl0iI
;
reg
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBo0iI
;
reg
[
TABITS
+
CORETSE_AHBlo1
:
0
]
CORETSE_AHBi0iI
;
wire
CORETSE_AHBO1iI
;
reg
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBI1iI
;
wire
CORETSE_AHBiOOI
;
reg
[
TABITS
:
0
]
CORETSE_AHBo1i
;
reg
CORETSE_AHBi1i
;
reg
CORETSE_AHBl1i
;
reg
CORETSE_AHBl1iI
;
reg
CORETSE_AHBI0oI
;
reg
CORETSE_AHBo1iI
;
reg
CORETSE_AHBi1iI
;
reg
CORETSE_AHBOoiI
;
reg
CORETSE_AHBIoiI
;
wire
CORETSE_AHBloiI
;
wire
CORETSE_AHBOIi
;
reg
CORETSE_AHBooiI
;
reg
CORETSE_AHBioiI
;
reg
CORETSE_AHBIIi
;
wire
CORETSE_AHBOOi
;
wire
CORETSE_AHBIOi
;
wire
CORETSE_AHBlOi
;
wire
CORETSE_AHBoOi
;
wire
CORETSE_AHBiOi
;
reg
CORETSE_AHBOiiI
;
reg
CORETSE_AHBIiiI
;
reg
CORETSE_AHBliiI
;
reg
[
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
:
0
]
CORETSE_AHBllOI
;
reg
CORETSE_AHBIlOI
;
reg
CORETSE_AHBoiiI
;
reg
CORETSE_AHBiiiI
;
reg
CORETSE_AHBOOOl
;
reg
CORETSE_AHBIOOl
;
wire
CORETSE_AHBlOOl
;
wire
CORETSE_AHBoOOl
;
//     generate logic as part of synthesis results.
wire
[
(
TABITS
-
1
)
:
0
]
#
1000
CORETSE_AHBoli
=
CORETSE_AHBO0iI
[
(
TABITS
+
(
CORETSE_AHBlo1
-
1
)
)
:
CORETSE_AHBlo1
]
;
assign
CORETSE_AHBlIiI
=
(
(
CORETSE_AHBIliI
[
(
TABITS
)
]
==
CORETSE_AHBlliI
[
(
TABITS
+
CORETSE_AHBlo1
)
]
)
&
(
CORETSE_AHBIliI
[
(
TABITS
-
1
)
:
0
]
>
CORETSE_AHBlliI
[
(
TABITS
+
CORETSE_AHBlo1
-
1
)
:
CORETSE_AHBlo1
]
)
)
|
(
(
CORETSE_AHBIliI
[
(
TABITS
)
]
!=
CORETSE_AHBlliI
[
(
TABITS
+
CORETSE_AHBlo1
)
]
)
&
(
CORETSE_AHBIliI
[
(
TABITS
-
1
)
:
0
]
<=
CORETSE_AHBlliI
[
(
TABITS
+
CORETSE_AHBlo1
-
1
)
:
CORETSE_AHBlo1
]
)
)
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBoIiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBoIiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIiI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBiIiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiIiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIiI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBOliI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
&
(
(
CORETSE_AHBolo
&
(
CORETSE_AHBo0iI
[
CORETSE_AHBlo1
-
1
:
0
]
==
{
CORETSE_AHBlo1
{
1
'h
1
}
}
)
)
|
CORETSE_AHBOIiI
[
1
]
|
CORETSE_AHBOIiI
[
5
]
|
CORETSE_AHBOIiI
[
3
]
)
)
CORETSE_AHBOliI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIiI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
else
if
(
CORETSE_AHBllo
)
case
(
CORETSE_AHBOIiI
)
6
'h
01
:
if
(
CORETSE_AHBoIiI
&
CORETSE_AHBOoiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
02
;
else
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
6
'h
02
:
if
(
CORETSE_AHBO0o
&
~
CORETSE_AHBIiiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
08
;
else
if
(
CORETSE_AHBolo
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
04
;
else
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
02
;
6
'h
04
:
if
(
~
CORETSE_AHBOliI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
08
;
else
if
(
CORETSE_AHBO0o
&
~
CORETSE_AHBIiiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
10
;
else
if
(
CORETSE_AHBilo
&
~
CORETSE_AHBOiiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
20
;
else
if
(
CORETSE_AHBOliI
&
~
CORETSE_AHBloiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
04
;
else
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
6
'h
08
:
if
(
CORETSE_AHBloiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
else
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
08
;
6
'h
10
:
if
(
~
CORETSE_AHBolo
&
~
CORETSE_AHBliiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
else
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
10
;
6
'h
20
:
if
(
CORETSE_AHBOliI
&
~
CORETSE_AHBloiI
)
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
20
;
else
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
default
:
CORETSE_AHBOIiI
<=
#
CORETSE_AHBIoII
6
'h
01
;
endcase
end
assign
CORETSE_AHBiOOI
=
CORETSE_AHBOoiI
|
~
CORETSE_AHBOIiI
[
0
]
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIIiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBIIiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIiI
[
1
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBOiiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBOiiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBilo
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIiiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBIiiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0o
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBliiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBliiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBolo
;
end
assign
CORETSE_AHBoliI
=
(
CORETSE_AHBiliI
[
(
TABITS
+
CORETSE_AHBlo1
)
:
0
]
+
1
)
;
assign
CORETSE_AHBo00I
=
(
{
CORETSE_AHBl0iI
[
(
TABITS
+
CORETSE_AHBlo1
)
:
CORETSE_AHBlo1
]
,
{
CORETSE_AHBlo1
{
1
'b
0
}
}
}
+
(
CORETSE_AHBIo1
/
8
)
)
;
assign
CORETSE_AHBl00I
=
(
CORETSE_AHBOIiI
[
4
]
)
?
CORETSE_AHBi0iI
:
(
(
CORETSE_AHBOIiI
[
2
]
|
CORETSE_AHBOIiI
[
3
]
|
CORETSE_AHBOIiI
[
5
]
)
&
CORETSE_AHBloiI
)
?
CORETSE_AHBo00I
:
(
CORETSE_AHBoIiI
&
(
(
(
|
CORETSE_AHBOIiI
[
2
:
1
]
)
&
CORETSE_AHBolo
)
|
CORETSE_AHBOIiI
[
3
]
|
CORETSE_AHBOIiI
[
5
]
)
)
?
CORETSE_AHBoliI
:
CORETSE_AHBiliI
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBiliI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiI
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBiliI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00I
;
end
assign
CORETSE_AHBlliI
=
CORETSE_AHBl00I
+
1
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBO0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiI
;
else
if
(
~
CORETSE_AHBlIII
[
TABITS
+
1
]
&
CORETSE_AHBlOOl
)
CORETSE_AHBO0iI
<=
#
CORETSE_AHBIoII
{
CORETSE_AHBlIII
[
TABITS
:
0
]
,
{
CORETSE_AHBlo1
{
1
'h
0
}
}
}
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBO0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBlliI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBI0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiI
;
else
CORETSE_AHBI0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0iI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBo0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiI
;
else
if
(
CORETSE_AHBllo
&
(
CORETSE_AHBolo
|
CORETSE_AHBOIiI
[
5
]
|
CORETSE_AHBOIiI
[
3
]
)
)
CORETSE_AHBo0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiliI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBi0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiI
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBOIiI
[
1
]
&
~
CORETSE_AHBIIiI
)
CORETSE_AHBi0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBl00I
;
end
assign
CORETSE_AHBO1iI
=
CORETSE_AHBiIiI
&
(
(
CORETSE_AHBolo
&
(
CORETSE_AHBo0iI
[
(
CORETSE_AHBlo1
-
1
)
:
0
]
==
{
CORETSE_AHBlo1
{
1
'h
1
}
}
)
)
|
CORETSE_AHBOIiI
[
1
]
|
CORETSE_AHBOIiI
[
5
]
|
CORETSE_AHBOIiI
[
3
]
)
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBI1iI
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
{
1
'b
0
}
}
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBO1iI
)
CORETSE_AHBI1iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBili
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBl0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBiOiI
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBO1iI
)
CORETSE_AHBl0iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0iI
;
end
assign
CORETSE_AHBiOi
=
CORETSE_AHBOIiI
[
1
]
;
assign
CORETSE_AHBloiI
=
CORETSE_AHBioiI
&
(
CORETSE_AHBooiI
|
(
CORETSE_AHBI1iI
[
CORETSE_AHBIo1
+
CORETSE_AHBlo1
]
&
(
CORETSE_AHBo0iI
[
(
CORETSE_AHBlo1
-
1
)
:
0
]
==
(
(
(
CORETSE_AHBIo1
/
8
)
-
1
)
-
CORETSE_AHBI1iI
[
CORETSE_AHBIo1
+:
CORETSE_AHBlo1
]
)
)
)
)
;
assign
CORETSE_AHBOIi
=
CORETSE_AHBloiI
&
~
CORETSE_AHBIIi
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIIi
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBIIi
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIiI
[
3
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBooiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
CORETSE_AHBooiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBloiI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBioiI
<=
#
CORETSE_AHBIoII
1
'b
1
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBooiI
)
CORETSE_AHBioiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBOIiI
[
2
]
)
CORETSE_AHBioiI
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
assign
CORETSE_AHBiio
=
CORETSE_AHBI1iI
[
CORETSE_AHBo0iI
[
(
CORETSE_AHBlo1
-
1
)
:
0
]
*
8
+:
8
]
;
assign
CORETSE_AHBOOi
=
CORETSE_AHBI1iI
[
CORETSE_AHBIo1
+
3
]
;
assign
CORETSE_AHBIOi
=
CORETSE_AHBI1iI
[
CORETSE_AHBIo1
+
4
]
;
assign
CORETSE_AHBlOi
=
CORETSE_AHBI1iI
[
CORETSE_AHBIo1
+
5
]
;
assign
CORETSE_AHBoOi
=
CORETSE_AHBI1iI
[
CORETSE_AHBIo1
+
7
]
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBi1i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
)
begin
if
(
CORETSE_AHBo1iI
)
CORETSE_AHBi1i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
(
~
CORETSE_AHBooiI
&
CORETSE_AHBloiI
)
|
(
~
CORETSE_AHBi1i
&
~
CORETSE_AHBo1iI
&
~
CORETSE_AHBI0o
&
(
CORETSE_AHBo1i
!=
CORETSE_AHBiliI
[
TABITS
+
CORETSE_AHBlo1
:
CORETSE_AHBlo1
]
)
)
)
CORETSE_AHBi1i
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBo1i
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBllo
&
~
CORETSE_AHBi1i
&
~
CORETSE_AHBo1iI
&
(
(
~
CORETSE_AHBooiI
&
CORETSE_AHBloiI
)
|
(
(
CORETSE_AHBo1i
!=
CORETSE_AHBiliI
[
TABITS
+
CORETSE_AHBlo1
:
CORETSE_AHBlo1
]
)
)
)
)
CORETSE_AHBo1i
<=
#
CORETSE_AHBIoII
CORETSE_AHBiliI
[
(
TABITS
+
CORETSE_AHBlo1
)
:
CORETSE_AHBlo1
]
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBl1i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
&
~
CORETSE_AHBl1iI
)
CORETSE_AHBl1i
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBl1iI
)
CORETSE_AHBl1i
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIliI
<=
#
CORETSE_AHBIoII
CORETSE_AHBol0I
;
else
if
(
CORETSE_AHBllo
&
CORETSE_AHBl1iI
&
~
CORETSE_AHBl1i
)
CORETSE_AHBIliI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOoi
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBi1iI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi1iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBloi
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBo1iI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo1iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBi1iI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBI0oI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI0oI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoi
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBl1iI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1iI
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0oI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBoiiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoiiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIII
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBiiiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiiiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBoiiI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBOOOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOOOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBiiiI
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIOOl
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIOOl
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOOl
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIlOI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIlOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIOOl
;
end
assign
CORETSE_AHBlOOl
=
CORETSE_AHBiiiI
&
~
CORETSE_AHBOOOl
;
assign
CORETSE_AHBoOOl
=
CORETSE_AHBIOOl
&
~
CORETSE_AHBIlOI
;
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBllOI
<=
#
CORETSE_AHBIoII
{
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
{
1
'b
0
}
}
;
else
if
(
~
CORETSE_AHBlIII
[
TABITS
+
1
]
&
CORETSE_AHBoOOl
)
CORETSE_AHBllOI
<=
#
CORETSE_AHBIoII
CORETSE_AHBili
;
else
if
(
CORETSE_AHBlIII
[
TABITS
+
1
]
&
CORETSE_AHBlOOl
)
CORETSE_AHBllOI
<=
#
CORETSE_AHBIoII
{
{
(
(
CORETSE_AHBIo1
+
CORETSE_AHBlo1
+
6
)
-
1
)
-
TABITS
{
1
'b
0
}
}
,
CORETSE_AHBlliI
[
TABITS
+
CORETSE_AHBlo1
:
CORETSE_AHBlo1
]
}
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBIoiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIoiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBOOII
;
end
always
@
(
posedge
CORETSE_AHBoi0
or
posedge
CORETSE_AHBO0II
)
begin
if
(
CORETSE_AHBO0II
)
CORETSE_AHBOoiI
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOoiI
<=
#
CORETSE_AHBIoII
CORETSE_AHBIoiI
;
end
endmodule
