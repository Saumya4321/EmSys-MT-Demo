// REVISION    : $Revision: 1.22 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2003, MENTOR
`timescale 1ns/1ns
module
pe_mcxmac
#
(
parameter
CORETSE_AHBlOI
=
1
'b
0
,
parameter
CORETSE_AHBiOI
=
1
'b
0
,
parameter
CORETSE_AHBoOI
=
1
'b
0
)
(
CORETSE_AHBO111
,
CORETSE_AHBI111
,
CORETSE_AHBl111
,
CORETSE_AHBiOO1
,
CORETSE_AHBoi0
,
CORETSE_AHBllo
,
CORETSE_AHBo111
,
CORETSE_AHBii0
,
CORETSE_AHBl0o
,
CORETSE_AHBol
,
CORETSE_AHBll
,
CORETSE_AHBo01
,
CORETSE_AHBiio
,
CORETSE_AHBiOi
,
CORETSE_AHBOIi
,
CORETSE_AHBIIi
,
CORETSE_AHBoOi
,
CORETSE_AHBlIi
,
CORETSE_AHBi111
,
CORETSE_AHBiIi
,
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
,
CORETSE_AHBI000
,
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
,
CORETSE_AHBiI
,
CORETSE_AHBlI
,
CORETSE_AHBIl
,
CORETSE_AHBoo01
,
CORETSE_AHBlOi
,
CORETSE_AHBOOi
,
CORETSE_AHBoo11
,
CORETSE_AHBIOi
,
CORETSE_AHBio1
,
CORETSE_AHBOi1
,
CORETSE_AHBIi1
,
CORETSE_AHBli1
,
CORETSE_AHBio11
,
CORETSE_AHBOi11
,
CORETSE_AHBoi1
,
CORETSE_AHBii1
,
CORETSE_AHBoo1
,
CORETSE_AHBll00
,
CORETSE_AHBIi11
,
CORETSE_AHBli11
,
CORETSE_AHBoi11
,
CORETSE_AHBii11
,
CORETSE_AHBoI
,
CORETSE_AHBII
,
CORETSE_AHBOl
,
CORETSE_AHBi01
,
CORETSE_AHBO11
,
CORETSE_AHBI11
,
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
,
CORETSE_AHBI0o
,
CORETSE_AHBIOo1
,
CORETSE_AHBlOo1
,
CORETSE_AHBoOo1
,
CORETSE_AHBIoo
,
CORETSE_AHBo0o
,
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
,
CORETSE_AHBiOo1
,
CORETSE_AHBOIo1
,
CORETSE_AHBo1o
,
CORETSE_AHBl1o
,
CORETSE_AHBIIo1
,
CORETSE_AHBlIo1
,
CORETSE_AHBiI00
,
CORETSE_AHBOl00
,
CORETSE_AHBIl00
,
CORETSE_AHBO1i
,
CORETSE_AHBI1i
,
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
,
CORETSE_AHBIlo1
,
CORETSE_AHBllo1
,
CORETSE_AHBolo1
,
CORETSE_AHBilo1
,
CORETSE_AHBO0o1
,
CORETSE_AHBI0o1
,
CORETSE_AHBl0o1
,
CORETSE_AHBo0o1
,
CORETSE_AHBi0o1
,
CORETSE_AHBO1o1
,
CORETSE_AHBI1o1
,
CORETSE_AHBl1o1
,
CORETSE_AHBo1o1
,
CORETSE_AHBi1o1
,
CORETSE_AHBOoo1
,
CORETSE_AHBIoo1
,
CORETSE_AHBloo1
,
CORETSE_AHBooo1
,
CORETSE_AHBioo1
,
CORETSE_AHBOio1
,
CORETSE_AHBIio1
,
CORETSE_AHBlio1
,
CORETSE_AHBoio1
,
CORETSE_AHBiio1
)
;
input
CORETSE_AHBO111
,
CORETSE_AHBI111
,
CORETSE_AHBl111
;
input
CORETSE_AHBiOO1
,
CORETSE_AHBoi0
,
CORETSE_AHBllo
;
input
CORETSE_AHBo111
,
CORETSE_AHBii0
,
CORETSE_AHBl0o
;
input
CORETSE_AHBol
,
CORETSE_AHBll
;
input
CORETSE_AHBo01
;
input
[
7
:
0
]
CORETSE_AHBiio
;
input
CORETSE_AHBiOi
,
CORETSE_AHBIIi
,
CORETSE_AHBOIi
;
input
CORETSE_AHBoOi
,
CORETSE_AHBlIi
;
input
[
15
:
0
]
CORETSE_AHBi111
;
input
CORETSE_AHBiIi
;
input
CORETSE_AHBI000
;
output
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
;
output
CORETSE_AHBOo11
,
CORETSE_AHBIo11
,
CORETSE_AHBlo11
;
output
[
1
:
0
]
CORETSE_AHBoo01
;
input
CORETSE_AHBiI
;
input
[
7
:
0
]
CORETSE_AHBlI
;
input
CORETSE_AHBIl
;
input
CORETSE_AHBlOi
,
CORETSE_AHBOOi
,
CORETSE_AHBoo11
,
CORETSE_AHBIOi
;
input
CORETSE_AHBio1
,
CORETSE_AHBOi1
,
CORETSE_AHBIi1
,
CORETSE_AHBli1
;
input
[
7
:
0
]
CORETSE_AHBoi1
;
input
[
31
:
0
]
CORETSE_AHBii1
;
input
CORETSE_AHBio11
;
input
[
4
:
0
]
CORETSE_AHBOi11
;
input
CORETSE_AHBoo1
;
output
[
47
:
0
]
CORETSE_AHBll00
;
output
CORETSE_AHBIi11
,
CORETSE_AHBli11
;
output
CORETSE_AHBoi11
,
CORETSE_AHBii11
;
output
CORETSE_AHBoI
;
output
[
7
:
0
]
CORETSE_AHBII
;
output
CORETSE_AHBOl
;
output
CORETSE_AHBi01
,
CORETSE_AHBO11
,
CORETSE_AHBI11
;
output
CORETSE_AHBolo
,
CORETSE_AHBOOo1
,
CORETSE_AHBO0o
,
CORETSE_AHBilo
;
output
CORETSE_AHBI0o
;
output
CORETSE_AHBIOo1
;
output
[
51
:
0
]
CORETSE_AHBlOo1
;
output
CORETSE_AHBoOo1
,
CORETSE_AHBIoo
;
output
[
7
:
0
]
CORETSE_AHBo0o
;
output
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
;
output
CORETSE_AHBiOo1
,
CORETSE_AHBOIo1
;
output
CORETSE_AHBo1o
;
output
[
32
:
0
]
CORETSE_AHBl1o
;
output
[
8
:
0
]
CORETSE_AHBIIo1
;
output
CORETSE_AHBlIo1
;
output
CORETSE_AHBiI00
,
CORETSE_AHBOl00
,
CORETSE_AHBIl00
;
output
[
31
:
0
]
CORETSE_AHBO1i
;
output
CORETSE_AHBI1i
;
output
CORETSE_AHBoIo1
,
CORETSE_AHBiIo1
,
CORETSE_AHBOlo1
;
output
CORETSE_AHBllo1
,
CORETSE_AHBolo1
,
CORETSE_AHBilo1
;
output
CORETSE_AHBIio1
,
CORETSE_AHBlio1
;
output
CORETSE_AHBoio1
,
CORETSE_AHBiio1
;
output
CORETSE_AHBIlo1
;
output
[
15
:
0
]
CORETSE_AHBO0o1
;
output
CORETSE_AHBI0o1
;
output
[
7
:
0
]
CORETSE_AHBl0o1
;
output
[
7
:
0
]
CORETSE_AHBo0o1
;
output
CORETSE_AHBi0o1
;
output
[
7
:
0
]
CORETSE_AHBO1o1
;
output
[
7
:
0
]
CORETSE_AHBI1o1
;
output
CORETSE_AHBl1o1
;
output
CORETSE_AHBo1o1
;
output
CORETSE_AHBi1o1
;
input
CORETSE_AHBOoo1
;
input
CORETSE_AHBIoo1
;
input
[
15
:
0
]
CORETSE_AHBloo1
;
input
CORETSE_AHBooo1
;
input
CORETSE_AHBOio1
;
input
[
79
:
0
]
CORETSE_AHBioo1
;
wire
CORETSE_AHBI0o1
;
wire
[
7
:
0
]
CORETSE_AHBl0o1
;
wire
[
7
:
0
]
CORETSE_AHBo0o1
;
wire
CORETSE_AHBi0o1
;
wire
[
7
:
0
]
CORETSE_AHBO1o1
;
wire
[
7
:
0
]
CORETSE_AHBI1o1
;
wire
CORETSE_AHBl1o1
;
wire
CORETSE_AHBo1o1
;
wire
CORETSE_AHBi1o1
;
wire
CORETSE_AHBOOi1
;
wire
CORETSE_AHBo1O1
;
wire
CORETSE_AHBi1O1
;
wire
CORETSE_AHBIOi1
,
CORETSE_AHBlOi1
;
wire
CORETSE_AHBoOi1
;
wire
CORETSE_AHBiOi1
;
wire
[
15
:
0
]
CORETSE_AHBOIi1
;
wire
CORETSE_AHBIIi1
,
CORETSE_AHBlIi1
;
wire
CORETSE_AHBoIi1
,
CORETSE_AHBiIi1
;
wire
[
47
:
0
]
CORETSE_AHBll00
;
wire
CORETSE_AHBOli1
,
CORETSE_AHBIli1
,
CORETSE_AHBlli1
;
wire
[
15
:
0
]
CORETSE_AHBoli1
;
wire
[
15
:
0
]
CORETSE_AHBili1
;
wire
[
15
:
0
]
CORETSE_AHBO0i1
;
wire
[
1
:
0
]
CORETSE_AHBoo01
,
CORETSE_AHBI0i1
;
wire
CORETSE_AHBl0i1
,
CORETSE_AHBo0i1
;
wire
CORETSE_AHBio01
,
CORETSE_AHBi0i1
,
CORETSE_AHBO1i1
;
wire
[
6
:
0
]
CORETSE_AHBI1i1
;
wire
[
6
:
0
]
CORETSE_AHBl1i1
,
CORETSE_AHBo1i1
;
wire
[
9
:
0
]
CORETSE_AHBi1i1
;
wire
[
3
:
0
]
CORETSE_AHBOoi1
;
wire
CORETSE_AHBIoi1
,
CORETSE_AHBloi1
;
wire
CORETSE_AHBooi1
,
CORETSE_AHBioi1
;
wire
[
15
:
0
]
CORETSE_AHBOii1
;
wire
[
7
:
0
]
CORETSE_AHBIii1
;
wire
[
3
:
0
]
CORETSE_AHBlii1
;
wire
[
3
:
0
]
CORETSE_AHBoii1
;
wire
CORETSE_AHBiii1
;
wire
CORETSE_AHBOOOo
,
CORETSE_AHBIOOo
;
wire
CORETSE_AHBiii0
,
CORETSE_AHBlOOo
;
wire
[
2
:
0
]
CORETSE_AHBoOOo
;
wire
CORETSE_AHBiOOo
,
CORETSE_AHBOIOo
;
wire
[
4
:
0
]
CORETSE_AHBIIOo
,
CORETSE_AHBlIOo
;
wire
CORETSE_AHBoIOo
;
wire
[
15
:
0
]
CORETSE_AHBiIOo
;
wire
CORETSE_AHBOlOo
,
CORETSE_AHBIlOo
;
wire
CORETSE_AHBllOo
,
CORETSE_AHBolOo
,
CORETSE_AHBilOo
,
CORETSE_AHBO0Oo
;
wire
CORETSE_AHBI0Oo
,
CORETSE_AHBl0Oo
;
wire
CORETSE_AHBIio1
,
CORETSE_AHBlio1
,
CORETSE_AHBo0Oo
,
CORETSE_AHBi0Oo
;
wire
CORETSE_AHBO1Oo
;
wire
CORETSE_AHBii01
;
assign
CORETSE_AHBO0o1
=
CORETSE_AHBOii1
;
assign
CORETSE_AHBili1
=
(
CORETSE_AHBO0i1
&
CORETSE_AHBi111
)
;
assign
CORETSE_AHBIlo1
=
CORETSE_AHBiii0
;
assign
CORETSE_AHBI0i1
=
{
(
CORETSE_AHBoo01
==
2
'b
10
)
,
(
CORETSE_AHBoo01
==
2
'b
00
|
CORETSE_AHBoo01
==
2
'b
01
)
}
;
assign
CORETSE_AHBI1Oo
=
CORETSE_AHBI1i1
;
pe_mcxmac_core
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
,
.CORETSE_AHBiOI
(
CORETSE_AHBiOI
)
,
.CORETSE_AHBlOI
(
CORETSE_AHBlOI
)
)
CORETSE_AHBl1Oo
(
.CORETSE_AHBiOO1
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBo1Oo
(
CORETSE_AHBllo
)
,
.CORETSE_AHBo111
(
CORETSE_AHBii0
)
,
.CORETSE_AHBi1Oo
(
CORETSE_AHBl0o
)
,
.CORETSE_AHBiI
(
CORETSE_AHBiI
)
,
.CORETSE_AHBlI
(
CORETSE_AHBlI
)
,
.CORETSE_AHBIl
(
CORETSE_AHBIl
)
,
.CORETSE_AHBol
(
CORETSE_AHBol
)
,
.CORETSE_AHBll
(
CORETSE_AHBll
)
,
.CORETSE_AHBiio
(
CORETSE_AHBiio
)
,
.CORETSE_AHBiOi
(
CORETSE_AHBiOi
)
,
.CORETSE_AHBIIi
(
CORETSE_AHBIIi
)
,
.CORETSE_AHBOIi
(
CORETSE_AHBOIi
)
,
.CORETSE_AHBlOi
(
CORETSE_AHBlOi
)
,
.CORETSE_AHBOOi
(
CORETSE_AHBOOi
)
,
.CORETSE_AHBoo11
(
CORETSE_AHBoo11
)
,
.CORETSE_AHBIOi
(
CORETSE_AHBIOi
)
,
.CORETSE_AHBoOi
(
CORETSE_AHBoOi
)
,
.CORETSE_AHBlIi
(
CORETSE_AHBlIi
)
,
.CORETSE_AHBi111
(
CORETSE_AHBili1
)
,
.CORETSE_AHBOoOo
(
CORETSE_AHBoli1
)
,
.CORETSE_AHBoo01
(
CORETSE_AHBI0i1
)
,
.CORETSE_AHBIOOo
(
CORETSE_AHBIOOo
)
,
.CORETSE_AHBOOOo
(
CORETSE_AHBOOOo
)
,
.CORETSE_AHBio01
(
CORETSE_AHBio01
)
,
.CORETSE_AHBoIi1
(
CORETSE_AHBoIi1
)
,
.CORETSE_AHBiIi1
(
CORETSE_AHBiIi1
)
,
.CORETSE_AHBll00
(
CORETSE_AHBll00
)
,
.CORETSE_AHBl0i1
(
CORETSE_AHBl0i1
)
,
.CORETSE_AHBo0i1
(
CORETSE_AHBo0i1
)
,
.CORETSE_AHBIoOo
(
CORETSE_AHBO1i1
)
,
.CORETSE_AHBlii1
(
CORETSE_AHBlii1
)
,
.CORETSE_AHBI1i1
(
CORETSE_AHBI1i1
)
,
.CORETSE_AHBl1i1
(
CORETSE_AHBl1i1
)
,
.CORETSE_AHBo1i1
(
CORETSE_AHBo1i1
)
,
.CORETSE_AHBi1i1
(
CORETSE_AHBi1i1
)
,
.CORETSE_AHBOoi1
(
CORETSE_AHBOoi1
)
,
.CORETSE_AHBoii1
(
CORETSE_AHBoii1
)
,
.CORETSE_AHBiii1
(
CORETSE_AHBiii1
)
,
.CORETSE_AHBIoi1
(
CORETSE_AHBIoi1
)
,
.CORETSE_AHBiIi
(
CORETSE_AHBooi1
)
,
.CORETSE_AHBioi1
(
CORETSE_AHBioi1
)
,
.CORETSE_AHBloOo
(
CORETSE_AHBOii1
)
,
.CORETSE_AHBi0i1
(
CORETSE_AHBi0i1
)
,
.CORETSE_AHBIii1
(
CORETSE_AHBIii1
)
,
.CORETSE_AHBloi1
(
CORETSE_AHBloi1
)
,
.CORETSE_AHBo0Oo
(
CORETSE_AHBo0Oo
)
,
.CORETSE_AHBi0Oo
(
CORETSE_AHBi0Oo
)
,
.CORETSE_AHBIio1
(
CORETSE_AHBIio1
)
,
.CORETSE_AHBlio1
(
CORETSE_AHBlio1
)
,
.CORETSE_AHBlli1
(
CORETSE_AHBlli1
)
,
.CORETSE_AHBlOOo
(
CORETSE_AHBlOOo
)
,
.CORETSE_AHBIli1
(
CORETSE_AHBIli1
)
,
.CORETSE_AHBiii0
(
CORETSE_AHBiii0
)
,
.CORETSE_AHBOli1
(
CORETSE_AHBOli1
)
,
.CORETSE_AHBolo
(
CORETSE_AHBolo
)
,
.CORETSE_AHBOOo1
(
CORETSE_AHBOOo1
)
,
.CORETSE_AHBO0o
(
CORETSE_AHBO0o
)
,
.CORETSE_AHBilo
(
CORETSE_AHBilo
)
,
.CORETSE_AHBI0o
(
CORETSE_AHBI0o
)
,
.CORETSE_AHBIoo
(
CORETSE_AHBIoo
)
,
.CORETSE_AHBoOo1
(
CORETSE_AHBoOo1
)
,
.CORETSE_AHBIOo1
(
CORETSE_AHBIOo1
)
,
.CORETSE_AHBlOo1
(
CORETSE_AHBlOo1
)
,
.CORETSE_AHBoOi1
(
CORETSE_AHBoOi1
)
,
.CORETSE_AHBoI
(
CORETSE_AHBoI
)
,
.CORETSE_AHBII
(
CORETSE_AHBII
)
,
.CORETSE_AHBOl
(
CORETSE_AHBOl
)
,
.CORETSE_AHBIOi1
(
CORETSE_AHBIOi1
)
,
.CORETSE_AHBlOi1
(
CORETSE_AHBlOi1
)
,
.CORETSE_AHBo0o
(
CORETSE_AHBo0o
)
,
.CORETSE_AHBi0o
(
CORETSE_AHBi0o
)
,
.CORETSE_AHBO1o
(
CORETSE_AHBO1o
)
,
.CORETSE_AHBI1o
(
CORETSE_AHBI1o
)
,
.CORETSE_AHBiOo1
(
CORETSE_AHBiOo1
)
,
.CORETSE_AHBOIo1
(
CORETSE_AHBOIo1
)
,
.CORETSE_AHBo1o
(
CORETSE_AHBo1o
)
,
.CORETSE_AHBl1o
(
CORETSE_AHBl1o
)
,
.CORETSE_AHBlIo1
(
CORETSE_AHBlIo1
)
,
.CORETSE_AHBIIo1
(
CORETSE_AHBIIo1
)
,
.CORETSE_AHBI0o1
(
CORETSE_AHBI0o1
)
,
.CORETSE_AHBl0o1
(
CORETSE_AHBl0o1
)
,
.CORETSE_AHBo0o1
(
CORETSE_AHBo0o1
)
,
.CORETSE_AHBi0o1
(
CORETSE_AHBi0o1
)
,
.CORETSE_AHBO1o1
(
CORETSE_AHBO1o1
)
,
.CORETSE_AHBI1o1
(
CORETSE_AHBI1o1
)
,
.CORETSE_AHBl1o1
(
CORETSE_AHBl1o1
)
,
.CORETSE_AHBo1o1
(
CORETSE_AHBo1o1
)
,
.CORETSE_AHBi1o1
(
CORETSE_AHBi1o1
)
,
.CORETSE_AHBOoo1
(
CORETSE_AHBOoo1
)
,
.CORETSE_AHBIoo1
(
CORETSE_AHBIoo1
)
,
.CORETSE_AHBloo1
(
CORETSE_AHBloo1
)
,
.CORETSE_AHBooo1
(
CORETSE_AHBooo1
)
,
.CORETSE_AHBOio1
(
CORETSE_AHBOio1
)
,
.CORETSE_AHBioo1
(
CORETSE_AHBioo1
)
,
.CORETSE_AHBiI00
(
CORETSE_AHBiI00
)
,
.CORETSE_AHBOl00
(
CORETSE_AHBOl00
)
,
.CORETSE_AHBIl00
(
CORETSE_AHBIl00
)
)
;
pemgt
CORETSE_AHBooOo
(
.CORETSE_AHBio11
(
CORETSE_AHBio11
)
,
.CORETSE_AHBoOOo
(
CORETSE_AHBoOOo
)
,
.CORETSE_AHBiOOo
(
CORETSE_AHBiOOo
)
,
.CORETSE_AHBOIOo
(
CORETSE_AHBOIOo
)
,
.CORETSE_AHBIIOo
(
CORETSE_AHBIIOo
)
,
.CORETSE_AHBlIOo
(
CORETSE_AHBlIOo
)
,
.CORETSE_AHBioOo
(
CORETSE_AHBoIOo
)
,
.CORETSE_AHBiIOo
(
CORETSE_AHBiIOo
)
,
.CORETSE_AHBOlOo
(
CORETSE_AHBOlOo
)
,
.CORETSE_AHBIlOo
(
CORETSE_AHBIlOo
)
,
.CORETSE_AHBo01
(
CORETSE_AHBo01
)
,
.CORETSE_AHBO1Oo
(
CORETSE_AHBO1Oo
)
,
.CORETSE_AHBi01
(
CORETSE_AHBi01
)
,
.CORETSE_AHBO11
(
CORETSE_AHBO11
)
,
.CORETSE_AHBI11
(
CORETSE_AHBI11
)
,
.CORETSE_AHBiOi1
(
CORETSE_AHBiOi1
)
,
.CORETSE_AHBOIi1
(
CORETSE_AHBOIi1
)
,
.CORETSE_AHBOiOo
(
)
,
.CORETSE_AHBIiOo
(
)
,
.CORETSE_AHBIIi1
(
CORETSE_AHBIIi1
)
,
.CORETSE_AHBlIi1
(
CORETSE_AHBlIi1
)
)
;
pehst
CORETSE_AHBliOo
(
.CORETSE_AHBio1
(
CORETSE_AHBio1
)
,
.CORETSE_AHBOi1
(
CORETSE_AHBOi1
)
,
.CORETSE_AHBIi1
(
CORETSE_AHBIi1
)
,
.CORETSE_AHBli1
(
CORETSE_AHBli1
)
,
.CORETSE_AHBoi1
(
CORETSE_AHBoi1
)
,
.CORETSE_AHBii1
(
CORETSE_AHBii1
)
,
.CORETSE_AHBOIi1
(
CORETSE_AHBOIi1
)
,
.CORETSE_AHBOi11
(
CORETSE_AHBOi11
)
,
.CORETSE_AHBiOi1
(
CORETSE_AHBiOi1
)
,
.CORETSE_AHBIIi1
(
CORETSE_AHBIIi1
)
,
.CORETSE_AHBlIi1
(
CORETSE_AHBlIi1
)
,
.CORETSE_AHBiIi
(
CORETSE_AHBiIi
)
,
.CORETSE_AHBIOi1
(
CORETSE_AHBIOi1
)
,
.CORETSE_AHBlOi1
(
CORETSE_AHBlOi1
)
,
.CORETSE_AHBoOi1
(
CORETSE_AHBoOi1
)
,
.CORETSE_AHBI000
(
CORETSE_AHBI000
)
,
.CORETSE_AHBol00
(
CORETSE_AHBol00
)
,
.CORETSE_AHBil00
(
CORETSE_AHBil00
)
,
.CORETSE_AHBO000
(
CORETSE_AHBO000
)
,
.CORETSE_AHBOo11
(
CORETSE_AHBOo11
)
,
.CORETSE_AHBIo11
(
CORETSE_AHBIo11
)
,
.CORETSE_AHBlo11
(
CORETSE_AHBlo11
)
,
.CORETSE_AHBO1i
(
CORETSE_AHBO1i
)
,
.CORETSE_AHBI1i
(
CORETSE_AHBI1i
)
,
.CORETSE_AHBoIi1
(
CORETSE_AHBoIi1
)
,
.CORETSE_AHBiIi1
(
CORETSE_AHBiIi1
)
,
.CORETSE_AHBll00
(
CORETSE_AHBll00
)
,
.CORETSE_AHBOoOo
(
CORETSE_AHBoli1
)
,
.CORETSE_AHBi111
(
CORETSE_AHBO0i1
)
,
.CORETSE_AHBl0i1
(
CORETSE_AHBl0i1
)
,
.CORETSE_AHBo0i1
(
CORETSE_AHBo0i1
)
,
.CORETSE_AHBio01
(
CORETSE_AHBio01
)
,
.CORETSE_AHBi0i1
(
CORETSE_AHBi0i1
)
,
.CORETSE_AHBO1i1
(
CORETSE_AHBO1i1
)
,
.CORETSE_AHBI1i1
(
CORETSE_AHBI1i1
)
,
.CORETSE_AHBIii1
(
CORETSE_AHBIii1
)
,
.CORETSE_AHBOii1
(
CORETSE_AHBOii1
)
,
.CORETSE_AHBl1i1
(
CORETSE_AHBl1i1
)
,
.CORETSE_AHBo1i1
(
CORETSE_AHBo1i1
)
,
.CORETSE_AHBi1i1
(
CORETSE_AHBi1i1
)
,
.CORETSE_AHBOoi1
(
CORETSE_AHBOoi1
)
,
.CORETSE_AHBIoi1
(
CORETSE_AHBIoi1
)
,
.CORETSE_AHBooi1
(
CORETSE_AHBooi1
)
,
.CORETSE_AHBioi1
(
CORETSE_AHBioi1
)
,
.CORETSE_AHBloi1
(
CORETSE_AHBloi1
)
,
.CORETSE_AHBoo01
(
CORETSE_AHBoo01
)
,
.CORETSE_AHBoiOo
(
)
,
.CORETSE_AHBOli1
(
CORETSE_AHBOli1
)
,
.CORETSE_AHBIli1
(
CORETSE_AHBIli1
)
,
.CORETSE_AHBlii1
(
CORETSE_AHBlii1
)
,
.CORETSE_AHBoii1
(
CORETSE_AHBoii1
)
,
.CORETSE_AHBiii1
(
CORETSE_AHBiii1
)
,
.CORETSE_AHBlli1
(
CORETSE_AHBlli1
)
,
.CORETSE_AHBOOOo
(
CORETSE_AHBOOOo
)
,
.CORETSE_AHBIOOo
(
CORETSE_AHBIOOo
)
,
.CORETSE_AHBiii0
(
CORETSE_AHBiii0
)
,
.CORETSE_AHBlOOo
(
CORETSE_AHBlOOo
)
,
.CORETSE_AHBoOOo
(
CORETSE_AHBoOOo
)
,
.CORETSE_AHBiOOo
(
CORETSE_AHBiOOo
)
,
.CORETSE_AHBOIOo
(
CORETSE_AHBOIOo
)
,
.CORETSE_AHBoIo1
(
CORETSE_AHBoIo1
)
,
.CORETSE_AHBiIo1
(
CORETSE_AHBiIo1
)
,
.CORETSE_AHBOlo1
(
CORETSE_AHBOlo1
)
,
.CORETSE_AHBIIOo
(
CORETSE_AHBIIOo
)
,
.CORETSE_AHBlIOo
(
CORETSE_AHBlIOo
)
,
.CORETSE_AHBoIOo
(
CORETSE_AHBoIOo
)
,
.CORETSE_AHBiIOo
(
CORETSE_AHBiIOo
)
,
.CORETSE_AHBOlOo
(
CORETSE_AHBOlOo
)
,
.CORETSE_AHBIlOo
(
CORETSE_AHBIlOo
)
,
.CORETSE_AHBii01
(
CORETSE_AHBii01
)
,
.CORETSE_AHBllOo
(
CORETSE_AHBllOo
)
,
.CORETSE_AHBolOo
(
CORETSE_AHBolOo
)
,
.CORETSE_AHBilOo
(
CORETSE_AHBilOo
)
,
.CORETSE_AHBO0Oo
(
CORETSE_AHBO0Oo
)
,
.CORETSE_AHBI0Oo
(
CORETSE_AHBI0Oo
)
,
.CORETSE_AHBiiOo
(
)
,
.CORETSE_AHBl0Oo
(
CORETSE_AHBl0Oo
)
,
.CORETSE_AHBOOIo
(
)
,
.CORETSE_AHBIOIo
(
)
)
;
pecar
CORETSE_AHBlOIo
(
.CORETSE_AHBO111
(
CORETSE_AHBO111
)
,
.CORETSE_AHBI111
(
CORETSE_AHBI111
)
,
.CORETSE_AHBl111
(
CORETSE_AHBl111
)
,
.CORETSE_AHBiOO1
(
CORETSE_AHBiOO1
)
,
.CORETSE_AHBo1Oo
(
1
'b
1
)
,
.CORETSE_AHBoi0
(
CORETSE_AHBoi0
)
,
.CORETSE_AHBllo
(
CORETSE_AHBllo
)
,
.CORETSE_AHBo111
(
CORETSE_AHBo111
)
,
.CORETSE_AHBi1Oo
(
1
'b
1
)
,
.CORETSE_AHBii0
(
CORETSE_AHBii0
)
,
.CORETSE_AHBl0o
(
CORETSE_AHBl0o
)
,
.CORETSE_AHBio11
(
CORETSE_AHBio11
)
,
.CORETSE_AHBoOIo
(
CORETSE_AHBIi11
)
,
.CORETSE_AHBiOIo
(
CORETSE_AHBli11
)
,
.CORETSE_AHBo011
(
CORETSE_AHBiii0
)
,
.CORETSE_AHBOi1
(
CORETSE_AHBOi1
)
,
.CORETSE_AHBio1
(
CORETSE_AHBio1
)
,
.CORETSE_AHBii01
(
CORETSE_AHBii01
)
,
.CORETSE_AHBllOo
(
CORETSE_AHBllOo
)
,
.CORETSE_AHBolOo
(
CORETSE_AHBolOo
)
,
.CORETSE_AHBilOo
(
CORETSE_AHBilOo
)
,
.CORETSE_AHBO0Oo
(
CORETSE_AHBO0Oo
)
,
.CORETSE_AHBI0Oo
(
CORETSE_AHBI0Oo
)
,
.CORETSE_AHBOIIo
(
1
'b
0
)
,
.CORETSE_AHBIIIo
(
1
'b
0
)
,
.CORETSE_AHBl0Oo
(
CORETSE_AHBl0Oo
)
,
.CORETSE_AHBOOIo
(
1
'b
0
)
,
.CORETSE_AHBIOIo
(
1
'b
0
)
,
.CORETSE_AHBoo1
(
CORETSE_AHBoo1
)
,
.CORETSE_AHBIi11
(
CORETSE_AHBIi11
)
,
.CORETSE_AHBli11
(
CORETSE_AHBli11
)
,
.CORETSE_AHBoi11
(
CORETSE_AHBoi11
)
,
.CORETSE_AHBii11
(
CORETSE_AHBii11
)
,
.CORETSE_AHBoio1
(
CORETSE_AHBoio1
)
,
.CORETSE_AHBiio1
(
CORETSE_AHBiio1
)
,
.CORETSE_AHBIio1
(
CORETSE_AHBIio1
)
,
.CORETSE_AHBlio1
(
CORETSE_AHBlio1
)
,
.CORETSE_AHBo0Oo
(
CORETSE_AHBo0Oo
)
,
.CORETSE_AHBi0Oo
(
CORETSE_AHBi0Oo
)
,
.CORETSE_AHBO1Oo
(
CORETSE_AHBO1Oo
)
,
.CORETSE_AHBII11
(
)
,
.CORETSE_AHBoI11
(
)
,
.CORETSE_AHBllo1
(
CORETSE_AHBllo1
)
,
.CORETSE_AHBolo1
(
CORETSE_AHBolo1
)
,
.CORETSE_AHBilo1
(
CORETSE_AHBilo1
)
,
.CORETSE_AHBlIIo
(
)
,
.CORETSE_AHBoIIo
(
)
,
.CORETSE_AHBiIIo
(
)
)
;
endmodule
