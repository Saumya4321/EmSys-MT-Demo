// REVISION    : $Revision: 1.1 $
//                   MENTOR Proprietary and Confidential
//                       Copyright (c) 2002, MENTOR
`timescale 1ps/1ps
module
mmcxwol
(
CORETSE_AHBii0
,
CORETSE_AHBl0o
,
CORETSE_AHBl0II
,
CORETSE_AHBo0o
,
CORETSE_AHBi0o
,
CORETSE_AHBO1o
,
CORETSE_AHBI1o
,
CORETSE_AHBl1o
,
CORETSE_AHBo1o
,
CORETSE_AHBiI00
,
CORETSE_AHBOl00
,
CORETSE_AHBIl00
,
CORETSE_AHBll00
,
CORETSE_AHBol00
,
CORETSE_AHBil00
,
CORETSE_AHBO000
,
CORETSE_AHBI000
)
;
input
CORETSE_AHBii0
;
input
CORETSE_AHBl0o
;
input
CORETSE_AHBl0II
;
input
[
7
:
0
]
CORETSE_AHBo0o
;
input
CORETSE_AHBi0o
;
input
CORETSE_AHBO1o
;
input
CORETSE_AHBI1o
;
input
[
22
:
20
]
CORETSE_AHBl1o
;
input
CORETSE_AHBo1o
;
input
CORETSE_AHBiI00
;
input
CORETSE_AHBOl00
;
input
CORETSE_AHBIl00
;
input
[
47
:
0
]
CORETSE_AHBll00
;
input
CORETSE_AHBol00
;
input
CORETSE_AHBil00
;
input
CORETSE_AHBO000
;
output
CORETSE_AHBI000
;
parameter
CORETSE_AHBIoII
=
1
;
reg
[
7
:
0
]
CORETSE_AHBl000
;
reg
[
7
:
0
]
CORETSE_AHBo000
;
reg
CORETSE_AHBli1I
;
reg
CORETSE_AHBoi1I
;
reg
CORETSE_AHBi000
;
reg
CORETSE_AHBO100
;
reg
CORETSE_AHBI100
;
reg
CORETSE_AHBii1I
;
reg
[
22
:
20
]
CORETSE_AHBl100
;
reg
CORETSE_AHBo100
;
reg
CORETSE_AHBi100
;
reg
CORETSE_AHBOo00
;
reg
CORETSE_AHBIo00
;
reg
CORETSE_AHBlo00
;
reg
[
3
:
0
]
CORETSE_AHBoo00
;
reg
[
4
:
0
]
CORETSE_AHBio00
;
reg
[
2
:
0
]
CORETSE_AHBOi00
;
reg
[
4
:
0
]
CORETSE_AHBIi00
;
wire
CORETSE_AHBli00
;
reg
CORETSE_AHBoi00
;
reg
CORETSE_AHBii00
;
wire
CORETSE_AHBOO10
;
reg
CORETSE_AHBIO10
;
reg
CORETSE_AHBlO10
;
reg
CORETSE_AHBI000
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl000
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBl000
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBli1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBli1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBi000
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBi000
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBO100
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBO100
<=
#
CORETSE_AHBIoII
CORETSE_AHBI1o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBl100
<=
#
CORETSE_AHBIoII
3
'b
000
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBl100
<=
#
CORETSE_AHBIoII
CORETSE_AHBl1o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBii1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBii1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBo1o
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBo100
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBo100
<=
#
CORETSE_AHBIoII
CORETSE_AHBiI00
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBi100
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBi100
<=
#
CORETSE_AHBIoII
CORETSE_AHBOl00
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOo00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBOo00
<=
#
CORETSE_AHBIoII
CORETSE_AHBIl00
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoi1I
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBoi1I
<=
#
CORETSE_AHBIoII
CORETSE_AHBli1I
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBo000
<=
#
CORETSE_AHBIoII
8
'h
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBo000
<=
#
CORETSE_AHBIoII
CORETSE_AHBl000
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBI100
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBI100
<=
#
CORETSE_AHBIoII
CORETSE_AHBO100
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIo00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBIo00
<=
#
CORETSE_AHBIoII
CORETSE_AHBO000
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBlo00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
)
CORETSE_AHBlo00
<=
#
CORETSE_AHBIoII
CORETSE_AHBIo00
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoo00
<=
#
CORETSE_AHBIoII
4
'd
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoi1I
&
CORETSE_AHBI100
)
CORETSE_AHBoo00
<=
#
CORETSE_AHBIoII
4
'd
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
CORETSE_AHBoo00
!=
4
'd
12
)
)
CORETSE_AHBoo00
<=
#
CORETSE_AHBIoII
CORETSE_AHBoo00
+
4
'd
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBio00
<=
#
CORETSE_AHBIoII
5
'd
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
(
CORETSE_AHBl000
!=
8
'h
FF
)
|
(
CORETSE_AHBoo00
!=
4
'd
12
)
|
CORETSE_AHBi000
)
)
CORETSE_AHBio00
<=
#
CORETSE_AHBIoII
5
'd
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
CORETSE_AHBl000
==
8
'h
FF
)
&
(
CORETSE_AHBoo00
==
4
'd
12
)
)
CORETSE_AHBio00
<=
#
CORETSE_AHBIoII
CORETSE_AHBio00
+
5
'd
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBOi00
<=
#
CORETSE_AHBIoII
3
'h
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
CORETSE_AHBi000
)
CORETSE_AHBOi00
<=
#
CORETSE_AHBIoII
3
'h
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
(
(
CORETSE_AHBio00
==
5
'd
6
)
&
(
CORETSE_AHBIi00
==
5
'h
0
)
)
|
(
CORETSE_AHBOi00
==
3
'h
6
)
)
)
CORETSE_AHBOi00
<=
#
CORETSE_AHBIoII
3
'h
1
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
CORETSE_AHBOi00
!=
3
'h
0
)
)
CORETSE_AHBOi00
<=
#
CORETSE_AHBIoII
CORETSE_AHBOi00
+
3
'h
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIi00
<=
#
CORETSE_AHBIoII
5
'h
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
CORETSE_AHBi000
)
CORETSE_AHBIi00
<=
#
CORETSE_AHBIoII
5
'h
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
(
(
CORETSE_AHBio00
==
5
'd
6
)
&
(
CORETSE_AHBIi00
==
5
'h
0
)
)
|
(
(
CORETSE_AHBOi00
==
3
'h
6
)
&
(
CORETSE_AHBIi00
==
5
'd
16
)
)
)
)
CORETSE_AHBIi00
<=
#
CORETSE_AHBIoII
5
'h
1
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBli1I
&
(
CORETSE_AHBOi00
==
3
'h
6
)
)
CORETSE_AHBIi00
<=
#
CORETSE_AHBIoII
CORETSE_AHBIi00
+
5
'h
1
;
end
assign
CORETSE_AHBli00
=
(
(
CORETSE_AHBOi00
==
3
'h
1
)
&
(
CORETSE_AHBll00
[
47
:
40
]
==
CORETSE_AHBo000
)
)
|
(
(
CORETSE_AHBOi00
==
3
'h
2
)
&
(
CORETSE_AHBll00
[
39
:
32
]
==
CORETSE_AHBo000
)
)
|
(
(
CORETSE_AHBOi00
==
3
'h
3
)
&
(
CORETSE_AHBll00
[
31
:
24
]
==
CORETSE_AHBo000
)
)
|
(
(
CORETSE_AHBOi00
==
3
'h
4
)
&
(
CORETSE_AHBll00
[
23
:
16
]
==
CORETSE_AHBo000
)
)
|
(
(
CORETSE_AHBOi00
==
3
'h
5
)
&
(
CORETSE_AHBll00
[
15
:
8
]
==
CORETSE_AHBo000
)
)
|
(
(
CORETSE_AHBOi00
==
3
'h
6
)
&
(
CORETSE_AHBll00
[
7
:
0
]
==
CORETSE_AHBo000
)
)
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBoi00
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoi1I
&
(
~
CORETSE_AHBli00
|
(
CORETSE_AHBOi00
==
3
'h
0
)
)
)
CORETSE_AHBoi00
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoi1I
&
CORETSE_AHBli00
&
CORETSE_AHBoi00
)
CORETSE_AHBoi00
<=
#
CORETSE_AHBIoII
1
'h
1
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBoi1I
&
CORETSE_AHBli00
&
(
CORETSE_AHBOi00
==
3
'h
1
)
&
(
CORETSE_AHBIi00
==
5
'd
1
)
)
CORETSE_AHBoi00
<=
#
CORETSE_AHBIoII
1
'h
1
;
end
assign
CORETSE_AHBOO10
=
(
CORETSE_AHBl0o
&
CORETSE_AHBli00
&
CORETSE_AHBoi00
&
(
CORETSE_AHBOi00
==
3
'h
6
)
&
(
CORETSE_AHBIi00
==
5
'd
16
)
)
;
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBii00
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
(
CORETSE_AHBoo00
==
4
'd
6
)
)
CORETSE_AHBii00
<=
#
CORETSE_AHBIoII
(
CORETSE_AHBOo00
|
CORETSE_AHBi100
|
CORETSE_AHBo100
)
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBIO10
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBii1I
)
CORETSE_AHBIO10
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBOO10
&
CORETSE_AHBii00
)
CORETSE_AHBIO10
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBlO10
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
(
CORETSE_AHBoo00
==
4
'd
6
)
)
CORETSE_AHBlO10
<=
#
CORETSE_AHBIoII
CORETSE_AHBOo00
;
end
always
@
(
posedge
CORETSE_AHBii0
or
posedge
CORETSE_AHBl0II
)
begin
if
(
CORETSE_AHBl0II
)
CORETSE_AHBI000
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBlo00
)
CORETSE_AHBI000
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
if
(
CORETSE_AHBl0o
&
CORETSE_AHBii1I
&
(
CORETSE_AHBl100
==
3
'b
000
)
&
(
(
CORETSE_AHBIO10
&
CORETSE_AHBil00
)
|
(
CORETSE_AHBlO10
&
CORETSE_AHBol00
)
)
)
CORETSE_AHBI000
<=
#
CORETSE_AHBIoII
1
'b
1
;
end
endmodule
