// REVISION    : $Revision: 1.22 $
//         Mentor Graphics Corporation Proprietary and Confidential
//         Copyright Mentor Graphics Corporation and Licensors 2004
module
mahbe_dual
#
(
parameter
CORETSE_AHBoOI
=
0
,
parameter
CORETSE_AHBOII
=
1
)
(
input
[
31
:
0
]
CORETSE_AHBloI0,
input
[
9
:
2
]
CORETSE_AHBooI0,
input
CORETSE_AHBioI0,
input
[
1
:
0
]
CORETSE_AHBOiI0,
input
CORETSE_AHBIiI0,
output
[
31
:
0
]
CORETSE_AHBliI0,
output
[
1
:
0
]
CORETSE_AHBoiI0,
output
CORETSE_AHBiiI0,
input
CORETSE_AHBOOl0,
input
CORETSE_AHBIOl0,
input
CORETSE_AHBlOl0,
input
[
1
:
0
]
CORETSE_AHBoOl0,
input
[
31
:
0
]
CORETSE_AHBiOl0,
output
CORETSE_AHBOIl0,
output
[
1
:
0
]
CORETSE_AHBIIl0,
output
[
31
:
2
]
CORETSE_AHBlIl0,
output
CORETSE_AHBoIl0,
output
[
31
:
0
]
CORETSE_AHBiIl0,
input
CORETSE_AHBOll0,
input
CORETSE_AHBIll0,
input
[
1
:
0
]
CORETSE_AHBlll0,
input
[
31
:
0
]
CORETSE_AHBoll0,
output
CORETSE_AHBill0,
output
[
1
:
0
]
CORETSE_AHBO0l0,
output
[
31
:
2
]
CORETSE_AHBI0l0,
output
CORETSE_AHBl0l0,
output
[
31
:
0
]
CORETSE_AHBo0l0,
input
CORETSE_AHBl1Il,
input
HCLK,
output
CORETSE_AHBiIll,
output
CORETSE_AHBOlll,
output
CORETSE_AHBIlll,
output
[
31
:
0
]
CORETSE_AHBllll,
output
[
1
:
0
]
CORETSE_AHBolll,
output
CORETSE_AHBilll,
output
CORETSE_AHBO0ll,
output
CORETSE_AHBI0ll,
output
[
1
:
0
]
CORETSE_AHBl0ll,
output
CORETSE_AHBo0ll,
input
CORETSE_AHBi0ll,
input
CORETSE_AHBO1ll,
input
CORETSE_AHBI1ll,
input
CORETSE_AHBl1ll,
input
CORETSE_AHBo1ll,
input
[
31
:
0
]
CORETSE_AHBi1ll,
input
[
1
:
0
]
CORETSE_AHBOoll,
output
CORETSE_AHBioOl,
output
CORETSE_AHBIoll,
output
[
7
:
0
]
CORETSE_AHBOiOl,
output
[
31
:
0
]
CORETSE_AHBloll,
input
[
31
:
0
]
CORETSE_AHBIiOl,
input
CORETSE_AHBliOl,
output
CORETSE_AHBi0l0,
input
CORETSE_AHBO1l0,
output
CORETSE_AHBooll,
output
[
5
:
0
]
CORETSE_AHBI1l0,
output
[
31
:
0
]
CORETSE_AHBl1l0,
output
[
31
:
0
]
CORETSE_AHBo1l0,
output
[
31
:
0
]
CORETSE_AHBi1l0,
output
[
31
:
0
]
CORETSE_AHBOol0,
output
[
31
:
0
]
CORETSE_AHBo00,
input
[
31
:
0
]
CORETSE_AHBl00,
input
[
15
:
0
]
CORETSE_AHBIIll,
input
[
31
:
0
]
CORETSE_AHBiIIl,
input
CORETSE_AHBOlIl,
output
CORETSE_AHBoIIl,
input
[
31
:
0
]
CORETSE_AHBllIl,
input
CORETSE_AHBolIl,
output
CORETSE_AHBIlIl,
input
[
31
:
0
]
CORETSE_AHBO0Il,
input
CORETSE_AHBI0Il,
output
CORETSE_AHBilIl
)
;
wire
[
31
:
0
]
CORETSE_AHBIol0
;
wire
CORETSE_AHBlol0
;
wire
CORETSE_AHBool0
;
wire
[
31
:
0
]
CORETSE_AHBlOIl
;
wire
CORETSE_AHBoOIl
;
wire
CORETSE_AHBIOIl
;
wire
[
31
:
0
]
CORETSE_AHBOIIl
;
wire
CORETSE_AHBIIIl
;
wire
CORETSE_AHBiOIl
;
wire
CORETSE_AHBlIIl
;
wire
[
31
:
0
]
CORETSE_AHBii0l
;
wire
[
31
:
0
]
CORETSE_AHBIO1l
;
dma_dual
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
,
.CORETSE_AHBOII
(
CORETSE_AHBOII
)
)
CORETSE_AHBiol0
(
.CORETSE_AHBl1Il
(
CORETSE_AHBl1Il
)
,
.HCLK
(
HCLK
)
,
.CORETSE_AHBo1Il
(
CORETSE_AHBIOl0
)
,
.CORETSE_AHBi1Il
(
CORETSE_AHBlOl0
)
,
.CORETSE_AHBOoIl
(
CORETSE_AHBoOl0
)
,
.CORETSE_AHBIoIl
(
CORETSE_AHBiOl0
)
,
.CORETSE_AHBloIl
(
CORETSE_AHBOIl0
)
,
.CORETSE_AHBooIl
(
CORETSE_AHBIIl0
)
,
.CORETSE_AHBioIl
(
CORETSE_AHBlIl0
)
,
.CORETSE_AHBOiIl
(
CORETSE_AHBoIl0
)
,
.CORETSE_AHBIiIl
(
CORETSE_AHBiIl0
)
,
.CORETSE_AHBIIll
(
CORETSE_AHBIIll
)
,
.CORETSE_AHBlIll
(
CORETSE_AHBii0l
)
,
.CORETSE_AHBoIll
(
CORETSE_AHBIO1l
)
,
.CORETSE_AHBliIl
(
CORETSE_AHBOll0
)
,
.CORETSE_AHBoiIl
(
CORETSE_AHBIll0
)
,
.CORETSE_AHBiiIl
(
CORETSE_AHBlll0
)
,
.CORETSE_AHBOOll
(
CORETSE_AHBoll0
)
,
.CORETSE_AHBIOll
(
CORETSE_AHBill0
)
,
.CORETSE_AHBlOll
(
CORETSE_AHBO0l0
)
,
.CORETSE_AHBoOll
(
CORETSE_AHBI0l0
)
,
.CORETSE_AHBiOll
(
CORETSE_AHBl0l0
)
,
.CORETSE_AHBOIll
(
CORETSE_AHBo0l0
)
,
.CORETSE_AHBiIll
(
CORETSE_AHBiIll
)
,
.CORETSE_AHBOlll
(
CORETSE_AHBOlll
)
,
.CORETSE_AHBIlll
(
CORETSE_AHBIlll
)
,
.CORETSE_AHBllll
(
CORETSE_AHBllll
)
,
.CORETSE_AHBolll
(
CORETSE_AHBolll
)
,
.CORETSE_AHBilll
(
CORETSE_AHBilll
)
,
.CORETSE_AHBi0ll
(
CORETSE_AHBi0ll
)
,
.CORETSE_AHBO1ll
(
CORETSE_AHBO1ll
)
,
.CORETSE_AHBI1ll
(
CORETSE_AHBI1ll
)
,
.CORETSE_AHBl1ll
(
CORETSE_AHBl1ll
)
,
.CORETSE_AHBo1ll
(
CORETSE_AHBo1ll
)
,
.CORETSE_AHBi1ll
(
CORETSE_AHBi1ll
)
,
.CORETSE_AHBOoll
(
CORETSE_AHBOoll
)
,
.CORETSE_AHBO0ll
(
CORETSE_AHBO0ll
)
,
.CORETSE_AHBI0ll
(
CORETSE_AHBI0ll
)
,
.CORETSE_AHBl0ll
(
CORETSE_AHBl0ll
)
,
.CORETSE_AHBo0ll
(
CORETSE_AHBo0ll
)
,
.CORETSE_AHBioOl
(
CORETSE_AHBIOIl
)
,
.CORETSE_AHBIoll
(
CORETSE_AHBIoll
)
,
.CORETSE_AHBOiOl
(
CORETSE_AHBOiOl
[
4
:
0
]
)
,
.CORETSE_AHBloll
(
CORETSE_AHBloll
)
,
.CORETSE_AHBIiOl
(
CORETSE_AHBlOIl
)
,
.CORETSE_AHBliOl
(
CORETSE_AHBoOIl
)
,
.CORETSE_AHBooll
(
CORETSE_AHBooll
)
)
;
slave
CORETSE_AHBOil0
(
.HWDATA
(
CORETSE_AHBloI0
)
,
.HADDR
(
CORETSE_AHBooI0
)
,
.HSEL
(
CORETSE_AHBioI0
)
,
.HTRANS
(
CORETSE_AHBOiI0
)
,
.HWRITE
(
CORETSE_AHBIiI0
)
,
.HCLK
(
HCLK
)
,
.CORETSE_AHBl1Il
(
CORETSE_AHBl1Il
)
,
.HREADY
(
CORETSE_AHBOOl0
)
,
.HRDATA
(
CORETSE_AHBliI0
)
,
.HRESP
(
CORETSE_AHBoiI0
)
,
.CORETSE_AHBIil0
(
CORETSE_AHBiiI0
)
,
.CORETSE_AHBioOl
(
CORETSE_AHBool0
)
,
.CORETSE_AHBIoll
(
CORETSE_AHBIoll
)
,
.CORETSE_AHBlIIl
(
CORETSE_AHBlIIl
)
,
.CORETSE_AHBOiOl
(
CORETSE_AHBOiOl
)
,
.CORETSE_AHBloll
(
CORETSE_AHBloll
)
,
.CORETSE_AHBIiOl
(
CORETSE_AHBIol0
)
,
.CORETSE_AHBliOl
(
CORETSE_AHBlol0
)
,
.CORETSE_AHBi0l0
(
CORETSE_AHBi0l0
)
,
.CORETSE_AHBO1l0
(
CORETSE_AHBO1l0
)
)
;
decoder
CORETSE_AHBlil0
(
.CORETSE_AHBlIIl
(
CORETSE_AHBlIIl
)
,
.CORETSE_AHBOiOl
(
CORETSE_AHBOiOl
[
7
:
3
]
)
,
.CORETSE_AHBioOl
(
CORETSE_AHBool0
)
,
.CORETSE_AHBIiOl
(
CORETSE_AHBIol0
)
,
.CORETSE_AHBliOl
(
CORETSE_AHBlol0
)
,
.CORETSE_AHBoiOl
(
CORETSE_AHBioOl
)
,
.CORETSE_AHBiiOl
(
CORETSE_AHBIiOl
)
,
.CORETSE_AHBOOIl
(
CORETSE_AHBliOl
)
,
.CORETSE_AHBIOIl
(
CORETSE_AHBIOIl
)
,
.CORETSE_AHBlOIl
(
CORETSE_AHBlOIl
)
,
.CORETSE_AHBoOIl
(
CORETSE_AHBoOIl
)
,
.CORETSE_AHBiOIl
(
CORETSE_AHBiOIl
)
,
.CORETSE_AHBOIIl
(
CORETSE_AHBOIIl
)
,
.CORETSE_AHBIIIl
(
CORETSE_AHBIIIl
)
,
.CORETSE_AHBoIIl
(
CORETSE_AHBoIIl
)
,
.CORETSE_AHBiIIl
(
CORETSE_AHBiIIl
)
,
.CORETSE_AHBOlIl
(
CORETSE_AHBOlIl
)
,
.CORETSE_AHBIlIl
(
CORETSE_AHBIlIl
)
,
.CORETSE_AHBllIl
(
CORETSE_AHBllIl
)
,
.CORETSE_AHBolIl
(
CORETSE_AHBolIl
)
,
.CORETSE_AHBilIl
(
CORETSE_AHBilIl
)
,
.CORETSE_AHBO0Il
(
CORETSE_AHBO0Il
)
,
.CORETSE_AHBI0Il
(
CORETSE_AHBI0Il
)
)
;
tsm_sysreg
#
(
.CORETSE_AHBOII
(
CORETSE_AHBOII
)
,
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
)
CORETSE_AHBoil0
(
.CORETSE_AHBiil0
(
HCLK
)
,
.CORETSE_AHBOO00
(
CORETSE_AHBl1Il
)
,
.CORETSE_AHBIO00
(
CORETSE_AHBiOIl
)
,
.CORETSE_AHBlO00
(
CORETSE_AHBIoll
)
,
.CORETSE_AHBoO00
(
CORETSE_AHBOiOl
[
4
:
0
]
)
,
.CORETSE_AHBiO00
(
CORETSE_AHBloll
)
,
.CORETSE_AHBl00
(
CORETSE_AHBl00
)
,
.CORETSE_AHBI1l0
(
CORETSE_AHBI1l0
)
,
.CORETSE_AHBl1l0
(
CORETSE_AHBl1l0
)
,
.CORETSE_AHBo1l0
(
CORETSE_AHBo1l0
)
,
.CORETSE_AHBi1l0
(
CORETSE_AHBi1l0
)
,
.CORETSE_AHBOol0
(
CORETSE_AHBOol0
)
,
.CORETSE_AHBo00
(
CORETSE_AHBo00
)
,
.CORETSE_AHBOI00
(
CORETSE_AHBii0l
)
,
.CORETSE_AHBII00
(
CORETSE_AHBIO1l
)
,
.CORETSE_AHBlI00
(
CORETSE_AHBOIIl
)
,
.CORETSE_AHBoI00
(
CORETSE_AHBIIIl
)
)
;
endmodule
