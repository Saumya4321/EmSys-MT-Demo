//                        Proprietary and Confidential 
// REVISION    : $Revision: 1.8 $ 
module
si_sal
(
input
CORETSE_AHBioOoI,
input
CORETSE_AHBOiOoI,
input
[
6
:
0
]
CORETSE_AHBIiOoI,
input
CORETSE_AHBliOoI,
input
CORETSE_AHBoiOoI,
input
CORETSE_AHBiiOoI,
input
CORETSE_AHBOOIoI,
input
CORETSE_AHBIOIoI,
input
[
5
:
0
]
CORETSE_AHBlOIoI,
input
[
31
:
0
]
CORETSE_AHBoOIoI,
input
[
31
:
0
]
CORETSE_AHBiOIoI,
input
[
31
:
0
]
CORETSE_AHBOIIoI,
input
[
31
:
0
]
CORETSE_AHBIIIoI,
output
CORETSE_AHBlIIoI,
output
CORETSE_AHBoIIoI
)
;
wire
[
7
:
0
]
CORETSE_AHBiIIoI
;
wire
CORETSE_AHBOlIoI
;
reg
CORETSE_AHBIlIoI
;
wire
CORETSE_AHBllIoI
;
reg
CORETSE_AHBolIoI
;
reg
CORETSE_AHBOoOi
;
wire
CORETSE_AHBilIoI
;
assign
CORETSE_AHBlIIoI
=
CORETSE_AHBOoOi
;
assign
CORETSE_AHBiIIoI
=
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBoOIoI
[
7
:
0
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBoOIoI
[
15
:
8
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBoOIoI
[
23
:
16
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBoOIoI
[
31
:
24
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBiOIoI
[
7
:
0
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBiOIoI
[
15
:
8
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBiOIoI
[
23
:
16
]
|
{
8
{
~
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBiOIoI
[
31
:
24
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBOIIoI
[
7
:
0
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBOIIoI
[
15
:
8
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBOIIoI
[
23
:
16
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
~
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBOIIoI
[
31
:
24
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBIIIoI
[
7
:
0
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
~
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBIIIoI
[
15
:
8
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
~
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBIIIoI
[
23
:
16
]
|
{
8
{
CORETSE_AHBIiOoI
[
6
]
&
CORETSE_AHBIiOoI
[
5
]
&
CORETSE_AHBIiOoI
[
4
]
&
CORETSE_AHBIiOoI
[
3
]
}
}
&
CORETSE_AHBIIIoI
[
31
:
24
]
;
assign
CORETSE_AHBOlIoI
=
(
(
~
CORETSE_AHBIiOoI
[
2
]
&
~
CORETSE_AHBIiOoI
[
1
]
&
~
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
0
]
)
|
(
(
~
CORETSE_AHBIiOoI
[
2
]
&
~
CORETSE_AHBIiOoI
[
1
]
&
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
1
]
)
|
(
(
~
CORETSE_AHBIiOoI
[
2
]
&
CORETSE_AHBIiOoI
[
1
]
&
~
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
2
]
)
|
(
(
~
CORETSE_AHBIiOoI
[
2
]
&
CORETSE_AHBIiOoI
[
1
]
&
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
3
]
)
|
(
(
CORETSE_AHBIiOoI
[
2
]
&
~
CORETSE_AHBIiOoI
[
1
]
&
~
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
4
]
)
|
(
(
CORETSE_AHBIiOoI
[
2
]
&
~
CORETSE_AHBIiOoI
[
1
]
&
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
5
]
)
|
(
(
CORETSE_AHBIiOoI
[
2
]
&
CORETSE_AHBIiOoI
[
1
]
&
~
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
6
]
)
|
(
(
CORETSE_AHBIiOoI
[
2
]
&
CORETSE_AHBIiOoI
[
1
]
&
CORETSE_AHBIiOoI
[
0
]
)
&
CORETSE_AHBiIIoI
[
7
]
)
;
always
@
(
posedge
CORETSE_AHBioOoI
or
negedge
CORETSE_AHBOiOoI
)
begin
if
(
!
CORETSE_AHBOiOoI
)
CORETSE_AHBIlIoI
<=
1
'b
0
;
else
if
(
CORETSE_AHBliOoI
)
CORETSE_AHBIlIoI
<=
CORETSE_AHBOlIoI
;
else
CORETSE_AHBIlIoI
<=
CORETSE_AHBIlIoI
;
end
assign
CORETSE_AHBO0IoI
=
(
CORETSE_AHBlOIoI
[
0
]
&
CORETSE_AHBOOIoI
)
|
(
CORETSE_AHBlOIoI
[
1
]
&
CORETSE_AHBiiOoI
)
|
(
CORETSE_AHBlOIoI
[
2
]
&
CORETSE_AHBoiOoI
)
|
(
CORETSE_AHBlOIoI
[
3
]
)
|
(
CORETSE_AHBlOIoI
[
4
]
&
CORETSE_AHBIlIoI
&
!
CORETSE_AHBiiOoI
&
!
CORETSE_AHBOOIoI
)
|
(
CORETSE_AHBlOIoI
[
5
]
&
CORETSE_AHBIlIoI
&
CORETSE_AHBiiOoI
&
!
CORETSE_AHBOOIoI
)
;
always
@
(
posedge
CORETSE_AHBioOoI
or
negedge
CORETSE_AHBOiOoI
)
begin
if
(
!
CORETSE_AHBOiOoI
)
begin
CORETSE_AHBolIoI
<=
1
'b
0
;
CORETSE_AHBOoOi
<=
1
'b
0
;
end
else
begin
CORETSE_AHBolIoI
<=
CORETSE_AHBllIoI
;
CORETSE_AHBOoOi
<=
CORETSE_AHBilIoI
;
end
end
assign
CORETSE_AHBllIoI
=
~
CORETSE_AHBO0IoI
;
assign
CORETSE_AHBoIIoI
=
CORETSE_AHBolIoI
;
assign
CORETSE_AHBilIoI
=
CORETSE_AHBIOIoI
&
CORETSE_AHBolIoI
|
~
CORETSE_AHBIOIoI
&
CORETSE_AHBOoOi
;
endmodule
