//               centralization improves synthesis and layout development 
// REVISION    : $Revision: 1.1 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
msgmii_clkrst
(
CORETSE_AHBIi0
,
CORETSE_AHBll1
,
CORETSE_AHBli0
,
CORETSE_AHBoi0
,
CORETSE_AHBii0
,
CORETSE_AHBlO1
,
CORETSE_AHBiO1
,
CORETSE_AHBoO10
,
CORETSE_AHBiO10
,
CORETSE_AHBOI10
,
CORETSE_AHBlI1
,
CORETSE_AHBoI1
,
CORETSE_AHBoO1
)
;
input
CORETSE_AHBIi0
;
input
CORETSE_AHBll1
;
input
CORETSE_AHBli0
;
input
CORETSE_AHBoi0
;
input
CORETSE_AHBii0
;
input
CORETSE_AHBlO1
;
input
CORETSE_AHBiO1
;
output
CORETSE_AHBoO10
;
output
CORETSE_AHBiO10
;
output
CORETSE_AHBOI10
;
output
CORETSE_AHBlI1
;
output
CORETSE_AHBoI1
;
output
CORETSE_AHBoO1
;
`define CORETSE_AHBIoII  \
# \
1
reg
CORETSE_AHBII10
;
reg
CORETSE_AHBlI10
;
reg
CORETSE_AHBoI10
;
reg
CORETSE_AHBiI10
;
reg
CORETSE_AHBOl10
;
reg
CORETSE_AHBIl10
;
reg
CORETSE_AHBll10
;
reg
CORETSE_AHBol10
;
reg
CORETSE_AHBil10
;
reg
CORETSE_AHBO010
;
reg
CORETSE_AHBI010
;
reg
CORETSE_AHBl010
;
wire
CORETSE_AHBo010
;
reg
CORETSE_AHBoO1
;
always
@
(
posedge
CORETSE_AHBli0
)
begin
CORETSE_AHBII10
<=
`CORETSE_AHBIoII
CORETSE_AHBIi0
;
end
always
@
(
posedge
CORETSE_AHBli0
)
begin
CORETSE_AHBlI10
<=
`CORETSE_AHBIoII
CORETSE_AHBII10
;
end
assign
CORETSE_AHBoO10
=
CORETSE_AHBll1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIi0
|
CORETSE_AHBlI10
)
;
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBOl10
<=
`CORETSE_AHBIoII
CORETSE_AHBIi0
;
end
always
@
(
posedge
CORETSE_AHBii0
)
begin
CORETSE_AHBIl10
<=
`CORETSE_AHBIoII
CORETSE_AHBOl10
;
end
assign
CORETSE_AHBOI10
=
CORETSE_AHBll1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIi0
|
CORETSE_AHBIl10
)
;
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBoI10
<=
`CORETSE_AHBIoII
CORETSE_AHBIi0
;
end
always
@
(
posedge
CORETSE_AHBoi0
)
begin
CORETSE_AHBiI10
<=
`CORETSE_AHBIoII
CORETSE_AHBoI10
;
end
assign
CORETSE_AHBiO10
=
CORETSE_AHBll1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIi0
|
CORETSE_AHBiI10
)
;
always
@
(
posedge
CORETSE_AHBlO1
)
begin
CORETSE_AHBll10
<=
`CORETSE_AHBIoII
CORETSE_AHBIi0
;
end
always
@
(
posedge
CORETSE_AHBlO1
)
begin
CORETSE_AHBol10
<=
`CORETSE_AHBIoII
CORETSE_AHBll10
;
end
assign
CORETSE_AHBlI1
=
CORETSE_AHBll1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIi0
|
CORETSE_AHBol10
)
;
always
@
(
posedge
CORETSE_AHBiO1
)
begin
CORETSE_AHBil10
<=
`CORETSE_AHBIoII
CORETSE_AHBIi0
;
end
always
@
(
posedge
CORETSE_AHBiO1
)
begin
CORETSE_AHBO010
<=
`CORETSE_AHBIoII
CORETSE_AHBil10
;
end
assign
CORETSE_AHBoI1
=
CORETSE_AHBll1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIi0
|
CORETSE_AHBO010
)
;
always
@
(
negedge
CORETSE_AHBiO1
)
begin
CORETSE_AHBI010
<=
`CORETSE_AHBIoII
CORETSE_AHBIi0
;
end
always
@
(
negedge
CORETSE_AHBiO1
)
begin
CORETSE_AHBl010
<=
`CORETSE_AHBIoII
CORETSE_AHBI010
;
end
assign
CORETSE_AHBo010
=
CORETSE_AHBll1
?
CORETSE_AHBIi0
:
(
CORETSE_AHBIi0
|
CORETSE_AHBl010
)
;
always
@
(
negedge
CORETSE_AHBiO1
or
posedge
CORETSE_AHBo010
)
begin
if
(
CORETSE_AHBo010
)
CORETSE_AHBoO1
<=
`CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoO1
<=
`CORETSE_AHBIoII
~
CORETSE_AHBoO1
;
end
endmodule
