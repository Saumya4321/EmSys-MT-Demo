//                        Proprietary and Confidential 
// REVISION    : $Revision: 1.7 $ 
module
tsm_sysreg
#
(
parameter
CORETSE_AHBOII
=
1
,
parameter
CORETSE_AHBoOI
=
0
)
(
input
CORETSE_AHBiil0,
input
CORETSE_AHBOO00,
input
CORETSE_AHBIO00,
input
CORETSE_AHBlO00,
input
[
4
:
0
]
CORETSE_AHBoO00,
input
[
31
:
0
]
CORETSE_AHBiO00,
input
[
31
:
0
]
CORETSE_AHBl00,
output
[
5
:
0
]
CORETSE_AHBI1l0,
output
[
31
:
0
]
CORETSE_AHBl1l0,
output
[
31
:
0
]
CORETSE_AHBo1l0,
output
[
31
:
0
]
CORETSE_AHBi1l0,
output
[
31
:
0
]
CORETSE_AHBOol0,
output
[
31
:
0
]
CORETSE_AHBo00,
output
[
31
:
0
]
CORETSE_AHBOI00,
output
[
31
:
0
]
CORETSE_AHBII00,
output
[
31
:
0
]
CORETSE_AHBlI00,
output
CORETSE_AHBoI00
)
;
wire
[
5
:
0
]
CORETSE_AHBoo0oI
;
wire
[
31
:
0
]
CORETSE_AHBio0oI
;
wire
[
31
:
0
]
CORETSE_AHBOi0oI
;
wire
[
31
:
0
]
CORETSE_AHBIi0oI
;
wire
[
31
:
0
]
CORETSE_AHBli0oI
;
wire
[
31
:
0
]
CORETSE_AHBoi0oI
;
reg
[
5
:
0
]
CORETSE_AHBii0oI
;
reg
[
31
:
0
]
CORETSE_AHBOO1oI
;
reg
[
31
:
0
]
CORETSE_AHBIO1oI
;
reg
[
31
:
0
]
CORETSE_AHBlO1oI
;
reg
[
31
:
0
]
CORETSE_AHBoO1oI
;
reg
[
31
:
0
]
CORETSE_AHBii
;
wire
CORETSE_AHBiO1oI
;
wire
CORETSE_AHBOI1oI
;
wire
[
31
:
0
]
CORETSE_AHBoi0l
;
reg
[
31
:
0
]
CORETSE_AHBii0l
;
wire
[
31
:
0
]
CORETSE_AHBOO1l
;
reg
[
31
:
0
]
CORETSE_AHBIO1l
;
`define CORETSE_AHBII1oI  \
5 \
'b \
1_0000
`define CORETSE_AHBlI1oI  \
5 \
'b \
1_0001
`define CORETSE_AHBoI1oI  \
5 \
'b \
1_0010
`define CORETSE_AHBiI1oI  \
5 \
'b \
1_0011
`define CORETSE_AHBOl1oI  \
5 \
'b \
1_0100
`define CORETSE_AHBIl1oI  \
5 \
'b \
1_0101
`define CORETSE_AHBll1oI  \
5 \
'b \
1_0110
`define CORETSE_AHBol1oI  \
5 \
'b \
1_1000
`define CORETSE_AHBil1oI  \
5 \
'b \
1_1001
assign
CORETSE_AHBI1l0
=
CORETSE_AHBii0oI
;
assign
CORETSE_AHBl1l0
=
CORETSE_AHBOO1oI
;
assign
CORETSE_AHBo1l0
=
CORETSE_AHBIO1oI
;
assign
CORETSE_AHBi1l0
=
CORETSE_AHBlO1oI
;
assign
CORETSE_AHBOol0
=
CORETSE_AHBoO1oI
;
assign
CORETSE_AHBo00
=
CORETSE_AHBii
;
generate
if
(
CORETSE_AHBOII
==
1
)
begin
assign
CORETSE_AHBOI00
=
CORETSE_AHBii0l
;
assign
CORETSE_AHBII00
=
CORETSE_AHBIO1l
;
end
else
begin
assign
CORETSE_AHBOI00
=
32
'b
0
;
assign
CORETSE_AHBII00
=
32
'b
0
;
end
endgenerate
assign
CORETSE_AHBO01oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBII1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBI01oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBlI1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBl01oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBoI1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBo01oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBiI1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBi01oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBOl1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBO11oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBIl1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBoo0oI
=
CORETSE_AHBO01oI
?
CORETSE_AHBiO00
[
5
:
0
]
:
CORETSE_AHBii0oI
;
assign
CORETSE_AHBio0oI
=
CORETSE_AHBI01oI
?
CORETSE_AHBiO00
:
CORETSE_AHBOO1oI
;
assign
CORETSE_AHBOi0oI
=
CORETSE_AHBl01oI
?
CORETSE_AHBiO00
:
CORETSE_AHBIO1oI
;
assign
CORETSE_AHBIi0oI
=
CORETSE_AHBo01oI
?
CORETSE_AHBiO00
:
CORETSE_AHBlO1oI
;
assign
CORETSE_AHBli0oI
=
CORETSE_AHBi01oI
?
CORETSE_AHBiO00
:
CORETSE_AHBoO1oI
;
assign
CORETSE_AHBoi0oI
=
CORETSE_AHBO11oI
?
CORETSE_AHBiO00
:
CORETSE_AHBii
;
generate
if
(
CORETSE_AHBOII
==
1
)
begin
assign
CORETSE_AHBiO1oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBol1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBOI1oI
=
(
!
CORETSE_AHBIO00
&&
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBil1oI
&&
!
CORETSE_AHBlO00
)
;
assign
CORETSE_AHBoi0l
=
CORETSE_AHBiO1oI
?
CORETSE_AHBiO00
:
CORETSE_AHBii0l
;
assign
CORETSE_AHBOO1l
=
CORETSE_AHBOI1oI
?
CORETSE_AHBiO00
:
CORETSE_AHBIO1l
;
end
endgenerate
generate
if
(
CORETSE_AHBOII
==
1
)
begin
assign
CORETSE_AHBoI00
=
CORETSE_AHBoO00
[
4
]
&&
(
!
(
&
CORETSE_AHBoO00
[
3
:
2
]
)
)
;
assign
CORETSE_AHBlI00
=
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBII1oI
)
}
}
&
{
26
'b
0
,
CORETSE_AHBii0oI
}
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBlI1oI
)
}
}
&
CORETSE_AHBOO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBoI1oI
)
}
}
&
CORETSE_AHBIO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBiI1oI
)
}
}
&
CORETSE_AHBlO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBOl1oI
)
}
}
&
CORETSE_AHBoO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBIl1oI
)
}
}
&
CORETSE_AHBii
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBll1oI
)
}
}
&
CORETSE_AHBl00
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBol1oI
)
}
}
&
CORETSE_AHBii0l
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBil1oI
)
}
}
&
CORETSE_AHBIO1l
)
;
end
else
begin
assign
CORETSE_AHBoI00
=
(
CORETSE_AHBoO00
[
4
:
3
]
==
2
'b
10
)
;
assign
CORETSE_AHBlI00
=
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBII1oI
)
}
}
&
{
26
'b
0
,
CORETSE_AHBii0oI
}
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBlI1oI
)
}
}
&
CORETSE_AHBOO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBoI1oI
)
}
}
&
CORETSE_AHBIO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBiI1oI
)
}
}
&
CORETSE_AHBlO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBOl1oI
)
}
}
&
CORETSE_AHBoO1oI
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBIl1oI
)
}
}
&
CORETSE_AHBii
)
|
(
{
32
{
(
CORETSE_AHBoO00
[
4
:
0
]
==
`CORETSE_AHBll1oI
)
}
}
&
CORETSE_AHBl00
)
;
end
endgenerate
generate
if
(
CORETSE_AHBOII
==
1
)
begin
always
@
(
posedge
CORETSE_AHBiil0
or
negedge
CORETSE_AHBOO00
)
begin
if
(
!
CORETSE_AHBOO00
)
begin
CORETSE_AHBii0l
<=
32
'h
FFFF_FFFF
;
CORETSE_AHBIO1l
<=
32
'h
FFFF_FFFF
;
end
else
begin
CORETSE_AHBii0l
<=
CORETSE_AHBoi0l
;
CORETSE_AHBIO1l
<=
CORETSE_AHBOO1l
;
end
end
end
endgenerate
always
@
(
posedge
CORETSE_AHBiil0
or
negedge
CORETSE_AHBOO00
)
begin
if
(
!
CORETSE_AHBOO00
)
begin
CORETSE_AHBii0oI
<=
6
'b
11_1111
;
CORETSE_AHBOO1oI
<=
32
'b
0
;
CORETSE_AHBIO1oI
<=
32
'b
0
;
CORETSE_AHBlO1oI
<=
32
'b
0
;
CORETSE_AHBoO1oI
<=
32
'b
0
;
CORETSE_AHBii
<=
32
'b
0
;
end
else
begin
CORETSE_AHBii0oI
<=
CORETSE_AHBoo0oI
;
CORETSE_AHBOO1oI
<=
CORETSE_AHBio0oI
;
CORETSE_AHBIO1oI
<=
CORETSE_AHBOi0oI
;
CORETSE_AHBlO1oI
<=
CORETSE_AHBIi0oI
;
CORETSE_AHBoO1oI
<=
CORETSE_AHBli0oI
;
CORETSE_AHBii
<=
CORETSE_AHBoi0oI
;
end
end
endmodule
