// REVISION    : $Revision: 1.13 $
//         Mentor Graphics Corporation Proprietary and Confidential
//         Copyright Mentor Graphics Corporation and Licensors 2004
`include "include.v"
module
dma_dual
#
(
parameter
CORETSE_AHBoOI
=
0
,
parameter
CORETSE_AHBOII
=
1
)
(
HCLK
,
CORETSE_AHBl1Il
,
CORETSE_AHBo1Il
,
CORETSE_AHBi1Il
,
CORETSE_AHBOoIl
,
CORETSE_AHBIoIl
,
CORETSE_AHBloIl
,
CORETSE_AHBooIl
,
CORETSE_AHBioIl
,
CORETSE_AHBOiIl
,
CORETSE_AHBIiIl
,
CORETSE_AHBliIl
,
CORETSE_AHBoiIl
,
CORETSE_AHBiiIl
,
CORETSE_AHBOOll
,
CORETSE_AHBIOll
,
CORETSE_AHBlOll
,
CORETSE_AHBoOll
,
CORETSE_AHBiOll
,
CORETSE_AHBOIll
,
CORETSE_AHBIIll
,
CORETSE_AHBlIll
,
CORETSE_AHBoIll
,
CORETSE_AHBiIll
,
CORETSE_AHBOlll
,
CORETSE_AHBIlll
,
CORETSE_AHBllll
,
CORETSE_AHBolll
,
CORETSE_AHBilll
,
CORETSE_AHBO0ll
,
CORETSE_AHBI0ll
,
CORETSE_AHBl0ll
,
CORETSE_AHBo0ll
,
CORETSE_AHBi0ll
,
CORETSE_AHBO1ll
,
CORETSE_AHBI1ll
,
CORETSE_AHBl1ll
,
CORETSE_AHBo1ll
,
CORETSE_AHBi1ll
,
CORETSE_AHBOoll
,
CORETSE_AHBioOl
,
CORETSE_AHBIoll
,
CORETSE_AHBOiOl
,
CORETSE_AHBloll
,
CORETSE_AHBIiOl
,
CORETSE_AHBliOl
,
CORETSE_AHBooll
)
;
input
CORETSE_AHBl1Il
;
input
HCLK
;
input
CORETSE_AHBo1Il
;
input
CORETSE_AHBi1Il
;
input
[
1
:
0
]
CORETSE_AHBOoIl
;
input
[
31
:
0
]
CORETSE_AHBIoIl
;
output
CORETSE_AHBloIl
;
output
[
1
:
0
]
CORETSE_AHBooIl
;
output
[
31
:
2
]
CORETSE_AHBioIl
;
output
CORETSE_AHBOiIl
;
output
[
31
:
0
]
CORETSE_AHBIiIl
;
input
CORETSE_AHBliIl
;
input
CORETSE_AHBoiIl
;
input
[
1
:
0
]
CORETSE_AHBiiIl
;
input
[
31
:
0
]
CORETSE_AHBOOll
;
output
CORETSE_AHBIOll
;
output
[
1
:
0
]
CORETSE_AHBlOll
;
output
[
31
:
2
]
CORETSE_AHBoOll
;
output
CORETSE_AHBiOll
;
output
[
31
:
0
]
CORETSE_AHBOIll
;
output
CORETSE_AHBiIll
;
output
CORETSE_AHBOlll
;
output
CORETSE_AHBIlll
;
output
[
31
:
0
]
CORETSE_AHBllll
;
output
[
1
:
0
]
CORETSE_AHBolll
;
input
CORETSE_AHBi0ll
;
output
CORETSE_AHBO0ll
;
output
CORETSE_AHBI0ll
;
output
[
1
:
0
]
CORETSE_AHBl0ll
;
output
CORETSE_AHBo0ll
;
output
CORETSE_AHBilll
;
input
CORETSE_AHBO1ll
;
input
CORETSE_AHBI1ll
;
input
CORETSE_AHBl1ll
;
input
CORETSE_AHBo1ll
;
input
[
31
:
0
]
CORETSE_AHBi1ll
;
input
[
1
:
0
]
CORETSE_AHBOoll
;
input
[
15
:
0
]
CORETSE_AHBIIll
;
input
CORETSE_AHBioOl
;
input
CORETSE_AHBIoll
;
input
[
4
:
0
]
CORETSE_AHBOiOl
;
input
[
31
:
0
]
CORETSE_AHBloll
;
output
[
31
:
0
]
CORETSE_AHBIiOl
;
output
CORETSE_AHBliOl
;
input
[
31
:
0
]
CORETSE_AHBlIll
;
input
[
31
:
0
]
CORETSE_AHBoIll
;
output
CORETSE_AHBooll
;
reg
CORETSE_AHBioll
;
reg
CORETSE_AHBOill
;
reg
CORETSE_AHBIill
;
reg
CORETSE_AHBlill
;
reg
CORETSE_AHBoill
;
reg
CORETSE_AHBiill
;
reg
CORETSE_AHBOO0l
;
reg
CORETSE_AHBIO0l
;
reg
CORETSE_AHBlO0l
;
reg
CORETSE_AHBoO0l
;
wire
CORETSE_AHBiO0l
;
wire
CORETSE_AHBOI0l
;
wire
CORETSE_AHBII0l
;
wire
CORETSE_AHBlI0l
;
reg
[
31
:
2
]
CORETSE_AHBoI0l
,
CORETSE_AHBiI0l
;
wire
[
31
:
2
]
CORETSE_AHBOl0l
,
CORETSE_AHBIl0l
;
reg
CORETSE_AHBll0l
;
wire
[
3
:
0
]
CORETSE_AHBol0l
;
wire
[
7
:
0
]
CORETSE_AHBil0l
;
wire
[
3
:
0
]
CORETSE_AHBO00l
;
wire
[
7
:
0
]
CORETSE_AHBI00l
;
reg
[
9
:
0
]
CORETSE_AHBl00l
;
reg
[
31
:
0
]
CORETSE_AHBIiOl
;
reg
CORETSE_AHBooll
;
wire
CORETSE_AHBo00l
,
CORETSE_AHBi00l
,
CORETSE_AHBO10l
;
wire
[
31
:
2
]
CORETSE_AHBI10l
;
wire
[
31
:
2
]
CORETSE_AHBl10l
;
wire
[
31
:
2
]
CORETSE_AHBo10l
,
CORETSE_AHBi10l
;
wire
CORETSE_AHBOo0l
;
wire
CORETSE_AHBIo0l
;
reg
CORETSE_AHBlo0l
;
reg
CORETSE_AHBoo0l
;
wire
[
7
:
0
]
CORETSE_AHBio0l
;
wire
[
7
:
0
]
CORETSE_AHBOi0l
;
reg
[
7
:
0
]
CORETSE_AHBIi0l
;
reg
[
7
:
0
]
CORETSE_AHBli0l
;
wire
[
31
:
0
]
CORETSE_AHBoi0l
;
reg
[
31
:
0
]
CORETSE_AHBii0l
;
wire
[
31
:
0
]
CORETSE_AHBOO1l
;
reg
[
31
:
0
]
CORETSE_AHBIO1l
;
generate
if
(
CORETSE_AHBOII
==
1
)
begin
assign
CORETSE_AHBoi0l
=
{
32
{
(
CORETSE_AHBii0l
==
CORETSE_AHBlIll
)
|
~
CORETSE_AHBl00l
[
8
]
}
}
&
32
'b
0
|
{
32
{
~
(
CORETSE_AHBii0l
==
CORETSE_AHBlIll
)
&
CORETSE_AHBl00l
[
8
]
}
}
&
(
CORETSE_AHBii0l
+
1
'b
1
)
;
assign
CORETSE_AHBOO1l
=
{
32
{
(
CORETSE_AHBIO1l
==
CORETSE_AHBoIll
)
|
~
CORETSE_AHBl00l
[
9
]
}
}
&
32
'b
0
|
{
32
{
~
(
CORETSE_AHBIO1l
==
CORETSE_AHBoIll
)
&
CORETSE_AHBl00l
[
9
]
}
}
&
(
CORETSE_AHBIO1l
+
1
'b
1
)
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBii0l
<=
32
'b
0
;
CORETSE_AHBIO1l
<=
32
'b
0
;
end
else
begin
CORETSE_AHBii0l
<=
CORETSE_AHBoi0l
;
CORETSE_AHBIO1l
<=
CORETSE_AHBOO1l
;
end
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
CORETSE_AHBlo0l
<=
1
'b
0
;
else
if
(
|
CORETSE_AHBil0l
==
1
'b
0
)
CORETSE_AHBlo0l
<=
1
'b
0
;
else
if
(
(
CORETSE_AHBil0l
==
CORETSE_AHBli0l
)
||
(
CORETSE_AHBii0l
==
CORETSE_AHBlIll
)
)
CORETSE_AHBlo0l
<=
1
'b
1
;
else
CORETSE_AHBlo0l
<=
CORETSE_AHBlo0l
;
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
CORETSE_AHBoo0l
<=
1
'b
0
;
else
if
(
|
CORETSE_AHBI00l
==
1
'b
0
)
CORETSE_AHBoo0l
<=
1
'b
0
;
else
if
(
(
CORETSE_AHBI00l
==
CORETSE_AHBIi0l
)
||
(
CORETSE_AHBIO1l
==
CORETSE_AHBoIll
)
)
CORETSE_AHBoo0l
<=
1
'b
1
;
else
CORETSE_AHBoo0l
<=
CORETSE_AHBoo0l
;
end
end
else
begin
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
CORETSE_AHBlo0l
<=
1
'b
0
;
else
if
(
|
CORETSE_AHBil0l
==
1
'b
0
)
CORETSE_AHBlo0l
<=
1
'b
0
;
else
if
(
CORETSE_AHBil0l
==
CORETSE_AHBli0l
)
CORETSE_AHBlo0l
<=
1
'b
1
;
else
CORETSE_AHBlo0l
<=
CORETSE_AHBlo0l
;
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
CORETSE_AHBoo0l
<=
1
'b
0
;
else
if
(
|
CORETSE_AHBI00l
==
1
'b
0
)
CORETSE_AHBoo0l
<=
1
'b
0
;
else
if
(
CORETSE_AHBI00l
==
CORETSE_AHBIi0l
)
CORETSE_AHBoo0l
<=
1
'b
1
;
else
CORETSE_AHBoo0l
<=
CORETSE_AHBoo0l
;
end
end
endgenerate
assign
CORETSE_AHBOi0l
=
(
!
CORETSE_AHBioOl
&&
~|
CORETSE_AHBOiOl
[
4
:
3
]
&&
!
CORETSE_AHBIoll
&&
CORETSE_AHBOiOl
[
2
:
0
]
==
`CORETSE_AHBlO1l
)
?
CORETSE_AHBloll
[
15
:
8
]
:
CORETSE_AHBli0l
;
assign
CORETSE_AHBio0l
=
(
!
CORETSE_AHBioOl
&&
~|
CORETSE_AHBOiOl
[
4
:
3
]
&&
!
CORETSE_AHBIoll
&&
CORETSE_AHBOiOl
[
2
:
0
]
==
`CORETSE_AHBoO1l
)
?
CORETSE_AHBloll
[
15
:
8
]
:
CORETSE_AHBIi0l
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBli0l
<=
8
'h
01
;
CORETSE_AHBIi0l
<=
8
'h
01
;
end
else
begin
CORETSE_AHBli0l
<=
CORETSE_AHBOi0l
;
CORETSE_AHBIi0l
<=
CORETSE_AHBio0l
;
end
end
assign
CORETSE_AHBO00l
=
{
CORETSE_AHBll0l
,
CORETSE_AHBoO0l
,
1
'b
0
,
|
CORETSE_AHBI00l
}
;
assign
CORETSE_AHBol0l
=
{
CORETSE_AHBll0l
,
1
'b
0
,
CORETSE_AHBlO0l
,
|
CORETSE_AHBil0l
}
;
always
@
(
*
)
begin
:
CORETSE_AHBiO1l
case
(
CORETSE_AHBOiOl
[
3
:
0
]
)
`CORETSE_AHBlO1l
:
CORETSE_AHBIiOl
=
{
16
'b
0
,
CORETSE_AHBli0l
,
7
'b
0
,
CORETSE_AHBII0l
}
;
`CORETSE_AHBOI1l
:
CORETSE_AHBIiOl
=
{
CORETSE_AHBoI0l
,
2
'b
0
}
;
`CORETSE_AHBII1l
:
CORETSE_AHBIiOl
=
{
8
'b
0
,
CORETSE_AHBil0l
,
12
'b
0
,
CORETSE_AHBol0l
}
;
`CORETSE_AHBoO1l
:
CORETSE_AHBIiOl
=
{
16
'b
0
,
CORETSE_AHBIi0l
,
7
'b
0
,
CORETSE_AHBlI0l
}
;
`CORETSE_AHBlI1l
:
CORETSE_AHBIiOl
=
{
CORETSE_AHBiI0l
,
2
'b
0
}
;
`CORETSE_AHBoI1l
:
CORETSE_AHBIiOl
=
{
8
'b
0
,
CORETSE_AHBI00l
,
12
'b
0
,
CORETSE_AHBO00l
}
;
`CORETSE_AHBiI1l
:
CORETSE_AHBIiOl
=
{
22
'b
0
,
CORETSE_AHBl00l
[
9
:
6
]
,
1
'b
0
,
CORETSE_AHBl00l
[
4
:
3
]
,
1
'b
0
,
CORETSE_AHBl00l
[
1
:
0
]
}
;
`CORETSE_AHBOl1l
:
CORETSE_AHBIiOl
=
{
22
'b
0
,
(
CORETSE_AHBl00l
&
{
CORETSE_AHBoo0l
,
CORETSE_AHBlo0l
,
CORETSE_AHBO00l
,
CORETSE_AHBol0l
}
)
}
;
default
:
CORETSE_AHBIiOl
=
32
'b
0
;
endcase
CORETSE_AHBooll
=
|
(
{
CORETSE_AHBl00l
[
9
:
8
]
,
CORETSE_AHBl00l
[
7
:
6
]
,
1
'b
0
,
CORETSE_AHBl00l
[
4
:
3
]
,
1
'b
0
,
CORETSE_AHBl00l
[
1
:
0
]
}
&
{
CORETSE_AHBoo0l
,
CORETSE_AHBlo0l
,
CORETSE_AHBO00l
,
CORETSE_AHBol0l
}
)
;
end
assign
CORETSE_AHBliOl
=
~
CORETSE_AHBOiOl
[
4
]
;
always
@
(
*
)
begin
:
CORETSE_AHBIl1l
CORETSE_AHBioll
=
0
;
CORETSE_AHBOill
=
0
;
CORETSE_AHBIill
=
0
;
CORETSE_AHBlill
=
0
;
CORETSE_AHBoill
=
0
;
CORETSE_AHBiill
=
0
;
CORETSE_AHBOO0l
=
0
;
CORETSE_AHBIO0l
=
0
;
if
(
!
CORETSE_AHBioOl
&&
~|
CORETSE_AHBOiOl
[
4
:
3
]
&&
!
CORETSE_AHBIoll
)
begin
case
(
CORETSE_AHBOiOl
[
2
:
0
]
)
`CORETSE_AHBlO1l
:
begin
CORETSE_AHBioll
=
CORETSE_AHBloll
[
0
]
;
CORETSE_AHBOill
=
!
CORETSE_AHBloll
[
0
]
;
end
`CORETSE_AHBOI1l
:
CORETSE_AHBoill
=
1
;
`CORETSE_AHBII1l
:
CORETSE_AHBOO0l
=
1
;
`CORETSE_AHBoO1l
:
begin
CORETSE_AHBIill
=
CORETSE_AHBloll
[
0
]
;
CORETSE_AHBlill
=
!
CORETSE_AHBloll
[
0
]
;
end
`CORETSE_AHBlI1l
:
CORETSE_AHBiill
=
1
;
`CORETSE_AHBoI1l
:
CORETSE_AHBIO0l
=
1
;
default
:
;
endcase
end
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
:
CORETSE_AHBll1l
if
(
!
CORETSE_AHBl1Il
)
CORETSE_AHBl00l
<=
0
;
else
if
(
!
CORETSE_AHBioOl
&&
~|
CORETSE_AHBOiOl
[
4
:
3
]
&&
CORETSE_AHBOiOl
[
2
:
0
]
==
`CORETSE_AHBiI1l
&&
!
CORETSE_AHBIoll
)
CORETSE_AHBl00l
<=
CORETSE_AHBloll
[
9
:
0
]
;
end
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
begin
CORETSE_AHBoI0l
<=
0
;
CORETSE_AHBiI0l
<=
0
;
CORETSE_AHBoO0l
<=
0
;
CORETSE_AHBlO0l
<=
0
;
end
else
begin
CORETSE_AHBoO0l
<=
CORETSE_AHBoO0l
&&
!
(
CORETSE_AHBIO0l
&&
CORETSE_AHBloll
[
2
]
)
||
CORETSE_AHBIo0l
;
CORETSE_AHBlO0l
<=
CORETSE_AHBlO0l
&&
!
(
CORETSE_AHBOO0l
&&
CORETSE_AHBloll
[
1
]
)
||
CORETSE_AHBOo0l
;
if
(
CORETSE_AHBoill
)
CORETSE_AHBoI0l
<=
CORETSE_AHBloll
[
31
:
2
]
;
else
CORETSE_AHBoI0l
<=
CORETSE_AHBo10l
;
if
(
CORETSE_AHBiill
)
CORETSE_AHBiI0l
<=
CORETSE_AHBloll
[
31
:
2
]
;
else
CORETSE_AHBiI0l
<=
CORETSE_AHBi10l
;
end
end
assign
CORETSE_AHBol1l
=
CORETSE_AHBOO0l
&&
CORETSE_AHBloll
[
0
]
;
assign
CORETSE_AHBil1l
=
CORETSE_AHBIO0l
&&
CORETSE_AHBloll
[
0
]
;
assign
CORETSE_AHBo00l
=
CORETSE_AHBi00l
||
CORETSE_AHBO10l
;
assign
CORETSE_AHBI10l
=
CORETSE_AHBoI0l
;
assign
CORETSE_AHBl10l
=
CORETSE_AHBiI0l
;
always
@
(
posedge
HCLK
or
negedge
CORETSE_AHBl1Il
)
begin
if
(
!
CORETSE_AHBl1Il
)
CORETSE_AHBll0l
<=
0
;
else
CORETSE_AHBll0l
<=
CORETSE_AHBll0l
&&
!
(
(
CORETSE_AHBOO0l
|
CORETSE_AHBIO0l
)
&&
CORETSE_AHBloll
[
3
]
)
||
CORETSE_AHBo00l
;
end
dmatx
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
)
CORETSE_AHBO01l
(
.CORETSE_AHBI01l
(
CORETSE_AHBo1Il
)
,
.HREADY
(
CORETSE_AHBi1Il
)
,
.HRESP
(
CORETSE_AHBOoIl
)
,
.HRDATA
(
CORETSE_AHBIoIl
)
,
.CORETSE_AHBl1Il
(
CORETSE_AHBl1Il
)
,
.HCLK
(
HCLK
)
,
.CORETSE_AHBl01l
(
CORETSE_AHBloIl
)
,
.HTRANS
(
CORETSE_AHBooIl
)
,
.HADDR
(
CORETSE_AHBioIl
)
,
.HWRITE
(
CORETSE_AHBOiIl
)
,
.HWDATA
(
CORETSE_AHBIiIl
)
,
.CORETSE_AHBi00l
(
CORETSE_AHBi00l
)
,
.CORETSE_AHBOo0l
(
CORETSE_AHBOo0l
)
,
.CORETSE_AHBo10l
(
CORETSE_AHBo10l
)
,
.CORETSE_AHBil0l
(
CORETSE_AHBil0l
)
,
.CORETSE_AHBioll
(
CORETSE_AHBioll
)
,
.CORETSE_AHBII0l
(
CORETSE_AHBII0l
)
,
.CORETSE_AHBOill
(
CORETSE_AHBOill
)
,
.CORETSE_AHBol1l
(
CORETSE_AHBol1l
)
,
.CORETSE_AHBI10l
(
CORETSE_AHBI10l
)
,
.CORETSE_AHBiIll
(
CORETSE_AHBiIll
)
,
.CORETSE_AHBOlll
(
CORETSE_AHBOlll
)
,
.CORETSE_AHBIlll
(
CORETSE_AHBIlll
)
,
.CORETSE_AHBllll
(
CORETSE_AHBllll
)
,
.CORETSE_AHBolll
(
CORETSE_AHBolll
)
,
.CORETSE_AHBO0ll
(
CORETSE_AHBO0ll
)
,
.CORETSE_AHBI0ll
(
CORETSE_AHBI0ll
)
,
.CORETSE_AHBl0ll
(
CORETSE_AHBl0ll
)
,
.CORETSE_AHBo0ll
(
CORETSE_AHBo0ll
)
,
.CORETSE_AHBi0ll
(
CORETSE_AHBi0ll
)
,
.CORETSE_AHBO1ll
(
CORETSE_AHBO1ll
)
)
;
dmarx
#
(
.CORETSE_AHBoOI
(
CORETSE_AHBoOI
)
)
CORETSE_AHBo01l
(
.CORETSE_AHBI01l
(
CORETSE_AHBliIl
)
,
.HREADY
(
CORETSE_AHBoiIl
)
,
.HRESP
(
CORETSE_AHBiiIl
)
,
.HRDATA
(
CORETSE_AHBOOll
)
,
.CORETSE_AHBl1Il
(
CORETSE_AHBl1Il
)
,
.HCLK
(
HCLK
)
,
.CORETSE_AHBl01l
(
CORETSE_AHBIOll
)
,
.HTRANS
(
CORETSE_AHBlOll
)
,
.HADDR
(
CORETSE_AHBoOll
)
,
.HWRITE
(
CORETSE_AHBiOll
)
,
.HWDATA
(
CORETSE_AHBOIll
)
,
.CORETSE_AHBO10l
(
CORETSE_AHBO10l
)
,
.CORETSE_AHBlI0l
(
CORETSE_AHBlI0l
)
,
.CORETSE_AHBIo0l
(
CORETSE_AHBIo0l
)
,
.CORETSE_AHBi10l
(
CORETSE_AHBi10l
)
,
.CORETSE_AHBI00l
(
CORETSE_AHBI00l
)
,
.CORETSE_AHBIill
(
CORETSE_AHBIill
)
,
.CORETSE_AHBlill
(
CORETSE_AHBlill
)
,
.CORETSE_AHBil1l
(
CORETSE_AHBil1l
)
,
.CORETSE_AHBl10l
(
CORETSE_AHBl10l
)
,
.CORETSE_AHBIIll
(
CORETSE_AHBIIll
)
,
.CORETSE_AHBilll
(
CORETSE_AHBilll
)
,
.CORETSE_AHBI1ll
(
CORETSE_AHBI1ll
)
,
.CORETSE_AHBl1ll
(
CORETSE_AHBl1ll
)
,
.CORETSE_AHBo1ll
(
CORETSE_AHBo1ll
)
,
.CORETSE_AHBi1ll
(
CORETSE_AHBi1ll
)
,
.CORETSE_AHBOoll
(
CORETSE_AHBOoll
)
)
;
endmodule
