// REVISION    : $Revision: 1.2 $
// Mentor Graphics Corporation Proprietary and Confidential
// Copyright 2007 Mentor Graphics Corporation and Licensors
`timescale 1ps/1ps
module
peanx_sync
(
CORETSE_AHBiOO1
,
CORETSE_AHBOo1
,
CORETSE_AHBOIO1
,
CORETSE_AHBIIO1
,
CORETSE_AHBlIO1
,
CORETSE_AHBiIO1
,
CORETSE_AHBOlO1
,
CORETSE_AHBllO1
,
CORETSE_AHBilO1
,
CORETSE_AHBO0O1
,
CORETSE_AHBI0O1
,
CORETSE_AHBl0O1
,
CORETSE_AHBo0O1
,
CORETSE_AHBi0O1
,
CORETSE_AHBO1O1
,
CORETSE_AHBI1O1
,
CORETSE_AHBOoI1
,
CORETSE_AHBloI1
,
CORETSE_AHBIoI1
,
CORETSE_AHBOiI1
,
CORETSE_AHBIiI1
,
CORETSE_AHBO0I1
,
CORETSE_AHBI0I1
,
CORETSE_AHBl0I1
,
CORETSE_AHBo1I1
,
CORETSE_AHBi1I1
,
CORETSE_AHBI1I1
,
CORETSE_AHBl1I1
,
CORETSE_AHBO1I1
,
CORETSE_AHBi0I1
,
CORETSE_AHBo101
,
CORETSE_AHBo0I1
)
;
input
CORETSE_AHBiOO1
;
input
CORETSE_AHBOo1
;
input
CORETSE_AHBOIO1
;
input
CORETSE_AHBIIO1
;
input
CORETSE_AHBlIO1
;
input
CORETSE_AHBiIO1
;
input
CORETSE_AHBOlO1
;
input
CORETSE_AHBllO1
;
input
CORETSE_AHBilO1
;
input
CORETSE_AHBO0O1
;
input
CORETSE_AHBI0O1
;
input
CORETSE_AHBl0O1
;
input
CORETSE_AHBo0O1
;
input
CORETSE_AHBi0O1
;
input
CORETSE_AHBO1O1
;
input
CORETSE_AHBI1O1
;
output
CORETSE_AHBOoI1
;
output
CORETSE_AHBIoI1
;
output
CORETSE_AHBloI1
;
output
CORETSE_AHBOiI1
;
output
CORETSE_AHBIiI1
;
output
CORETSE_AHBO0I1
;
output
CORETSE_AHBI0I1
;
output
CORETSE_AHBl0I1
;
output
CORETSE_AHBo1I1
;
output
CORETSE_AHBi1I1
;
output
CORETSE_AHBI1I1
;
output
CORETSE_AHBl1I1
;
output
CORETSE_AHBO1I1
;
output
CORETSE_AHBi0I1
;
output
CORETSE_AHBo101
;
output
CORETSE_AHBo0I1
;
reg
CORETSE_AHBOoI1
;
reg
CORETSE_AHBIoI1
;
reg
CORETSE_AHBloI1
;
reg
CORETSE_AHBOiI1
;
reg
CORETSE_AHBIiI1
;
reg
CORETSE_AHBO0I1
;
reg
CORETSE_AHBI0I1
;
reg
CORETSE_AHBl0I1
;
reg
CORETSE_AHBo1I1
;
reg
CORETSE_AHBi1I1
;
reg
CORETSE_AHBI1I1
;
reg
CORETSE_AHBl1I1
;
reg
CORETSE_AHBO1I1
;
reg
CORETSE_AHBi0I1
;
reg
CORETSE_AHBo101
;
reg
CORETSE_AHBo0I1
;
parameter
CORETSE_AHBIoII
=
1
;
reg
CORETSE_AHBOIlo
;
reg
CORETSE_AHBIIlo
;
reg
CORETSE_AHBlIlo
;
reg
CORETSE_AHBoIlo
;
reg
CORETSE_AHBiIlo
;
reg
CORETSE_AHBOllo
;
reg
CORETSE_AHBIllo
;
reg
CORETSE_AHBlllo
;
reg
CORETSE_AHBollo
;
reg
CORETSE_AHBillo
;
reg
CORETSE_AHBO0lo
;
reg
CORETSE_AHBI0lo
;
reg
CORETSE_AHBl0lo
;
reg
CORETSE_AHBo0lo
;
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOIlo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOIlo
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBO0I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO0I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIlo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBI0I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI0I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0I1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIIlo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIIlo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOlO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl0I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl0I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIlo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBlIlo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlIlo
<=
#
CORETSE_AHBIoII
CORETSE_AHBi0O1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo0I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo0I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIlo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBoIlo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBoIlo
<=
#
CORETSE_AHBIoII
CORETSE_AHBO1O1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo101
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBo101
<=
#
CORETSE_AHBIoII
CORETSE_AHBoIlo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBiIlo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBiIlo
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0O1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBi0I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBi0I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBiIlo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOllo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBOllo
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0O1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBO1I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBO1I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOllo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIllo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBIllo
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0O1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBI1I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBI1I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBIllo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBlllo
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBlllo
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0O1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl1I1
<=
#
CORETSE_AHBIoII
1
'b
0
;
else
CORETSE_AHBl1I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBlllo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBollo
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBollo
<=
#
CORETSE_AHBIoII
CORETSE_AHBllO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo1I1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBo1I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBollo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBillo
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBillo
<=
#
CORETSE_AHBIoII
CORETSE_AHBilO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBi1I1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBi1I1
<=
#
CORETSE_AHBIoII
CORETSE_AHBillo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBO0lo
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBO0lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOo1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOoI1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOoI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBO0lo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBI0lo
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBI0lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBOIO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIoI1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBIoI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBI0lo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBl0lo
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBl0lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBIIO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBloI1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBloI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBl0lo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBo0lo
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBo0lo
<=
#
CORETSE_AHBIoII
CORETSE_AHBlIO1
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBOiI1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBOiI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBo0lo
;
end
always
@
(
posedge
CORETSE_AHBiOO1
or
posedge
CORETSE_AHBI1O1
)
begin
if
(
CORETSE_AHBI1O1
)
CORETSE_AHBIiI1
<=
#
CORETSE_AHBIoII
1
'h
0
;
else
CORETSE_AHBIiI1
<=
#
CORETSE_AHBIoII
CORETSE_AHBOiI1
;
end
endmodule
